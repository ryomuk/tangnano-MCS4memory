//-----------------------------------------------------------------------------
//
// ROM image
//
//-----------------------------------------------------------------------------
module rom_image( addr, dout );
//-----------------------------------------------------------------------------
  input [11:0] addr;
  output [7:0] dout;
//-----------------------------------------------------------------------------
  reg [7:0]    rom [4095:0];
//-----------------------------------------------------------------------------
  assign dout = rom[addr];
  initial
    begin
    rom['h000]=8'hF0; rom['h001]=8'hD0; rom['h002]=8'hFD; rom['h003]=8'h59;
    rom['h004]=8'h39; rom['h005]=8'h5D; rom['h006]=8'h82; rom['h007]=8'h22;
    rom['h008]=8'h00; rom['h009]=8'hA3; rom['h00A]=8'h58; rom['h00B]=8'hEE;
    rom['h00C]=8'h58; rom['h00D]=8'hE2; rom['h00E]=8'h73; rom['h00F]=8'h09;
    rom['h010]=8'hF0; rom['h011]=8'h58; rom['h012]=8'hEE; rom['h013]=8'h20;
    rom['h014]=8'h3B; rom['h015]=8'h5E; rom['h016]=8'h00; rom['h017]=8'h20;
    rom['h018]=8'h17; rom['h019]=8'h5E; rom['h01A]=8'h00; rom['h01B]=8'h22;
    rom['h01C]=8'h5D; rom['h01D]=8'h5D; rom['h01E]=8'h28; rom['h01F]=8'h5D;
    rom['h020]=8'h00; rom['h021]=8'h5D; rom['h022]=8'h71; rom['h023]=8'h5C;
    rom['h024]=8'hEF; rom['h025]=8'h14; rom['h026]=8'h2B; rom['h027]=8'h5D;
    rom['h028]=8'h5C; rom['h029]=8'h40; rom['h02A]=8'h1B; rom['h02B]=8'h5D;
    rom['h02C]=8'h28; rom['h02D]=8'h20; rom['h02E]=8'h72; rom['h02F]=8'h5D;
    rom['h030]=8'hC3; rom['h031]=8'h1C; rom['h032]=8'h37; rom['h033]=8'h50;
    rom['h034]=8'h87; rom['h035]=8'h4C; rom['h036]=8'h06; rom['h037]=8'h20;
    rom['h038]=8'h77; rom['h039]=8'h5D; rom['h03A]=8'hC3; rom['h03B]=8'h1C;
    rom['h03C]=8'h41; rom['h03D]=8'h50; rom['h03E]=8'h87; rom['h03F]=8'h4C;
    rom['h040]=8'h30; rom['h041]=8'h20; rom['h042]=8'h52; rom['h043]=8'h5D;
    rom['h044]=8'hC3; rom['h045]=8'h1C; rom['h046]=8'h49; rom['h047]=8'h4C;
    rom['h048]=8'hAE; rom['h049]=8'h20; rom['h04A]=8'h57; rom['h04B]=8'h5D;
    rom['h04C]=8'hC3; rom['h04D]=8'h1C; rom['h04E]=8'h51; rom['h04F]=8'h4C;
    rom['h050]=8'h73; rom['h051]=8'h20; rom['h052]=8'h43; rom['h053]=8'h5D;
    rom['h054]=8'hC3; rom['h055]=8'h1C; rom['h056]=8'h59; rom['h057]=8'h4C;
    rom['h058]=8'hD5; rom['h059]=8'h20; rom['h05A]=8'h42; rom['h05B]=8'h5D;
    rom['h05C]=8'hC3; rom['h05D]=8'h1C; rom['h05E]=8'h61; rom['h05F]=8'h48;
    rom['h060]=8'hF3; rom['h061]=8'h20; rom['h062]=8'h67; rom['h063]=8'h5D;
    rom['h064]=8'hC3; rom['h065]=8'h1C; rom['h066]=8'h69; rom['h067]=8'h4C;
    rom['h068]=8'h00; rom['h069]=8'h20; rom['h06A]=8'h76; rom['h06B]=8'h5D;
    rom['h06C]=8'hC3; rom['h06D]=8'h1C; rom['h06E]=8'h71; rom['h06F]=8'h41;
    rom['h070]=8'h00; rom['h071]=8'h20; rom['h072]=8'h6C; rom['h073]=8'h5D;
    rom['h074]=8'hC3; rom['h075]=8'h1C; rom['h076]=8'h79; rom['h077]=8'h4A;
    rom['h078]=8'hD3; rom['h079]=8'h20; rom['h07A]=8'h4C; rom['h07B]=8'h5D;
    rom['h07C]=8'hC3; rom['h07D]=8'h1C; rom['h07E]=8'h81; rom['h07F]=8'h4B;
    rom['h080]=8'h1C; rom['h081]=8'h20; rom['h082]=8'h91; rom['h083]=8'h5E;
    rom['h084]=8'h00; rom['h085]=8'h40; rom['h086]=8'h1B; rom['h087]=8'h20;
    rom['h088]=8'h40; rom['h089]=8'h5E; rom['h08A]=8'h00; rom['h08B]=8'h5D;
    rom['h08C]=8'h00; rom['h08D]=8'h5D; rom['h08E]=8'h28; rom['h08F]=8'h5D;
    rom['h090]=8'hB7; rom['h091]=8'hA3; rom['h092]=8'hBA; rom['h093]=8'h20;
    rom['h094]=8'h47; rom['h095]=8'h5E; rom['h096]=8'h00; rom['h097]=8'h5D;
    rom['h098]=8'h00; rom['h099]=8'h5D; rom['h09A]=8'h28; rom['h09B]=8'h5D;
    rom['h09C]=8'hB7; rom['h09D]=8'hA3; rom['h09E]=8'hF1; rom['h09F]=8'hF5;
    rom['h0A0]=8'hF1; rom['h0A1]=8'hF5; rom['h0A2]=8'hBB; rom['h0A3]=8'h5D;
    rom['h0A4]=8'h5C; rom['h0A5]=8'hC0; rom['h0A6]=8'h2E; rom['h0A7]=8'h30;
    rom['h0A8]=8'h5D; rom['h0A9]=8'hD0; rom['h0AA]=8'h12; rom['h0AB]=8'hAD;
    rom['h0AC]=8'hC0; rom['h0AD]=8'h2E; rom['h0AE]=8'h3A; rom['h0AF]=8'h5D;
    rom['h0B0]=8'hD0; rom['h0B1]=8'h12; rom['h0B2]=8'hB4; rom['h0B3]=8'hC1;
    rom['h0B4]=8'h2E; rom['h0B5]=8'h41; rom['h0B6]=8'h5D; rom['h0B7]=8'hD0;
    rom['h0B8]=8'h12; rom['h0B9]=8'hBB; rom['h0BA]=8'hC0; rom['h0BB]=8'h2E;
    rom['h0BC]=8'h47; rom['h0BD]=8'h5D; rom['h0BE]=8'hD0; rom['h0BF]=8'h12;
    rom['h0C0]=8'hC2; rom['h0C1]=8'hC1; rom['h0C2]=8'h2E; rom['h0C3]=8'h61;
    rom['h0C4]=8'h5D; rom['h0C5]=8'hD0; rom['h0C6]=8'h12; rom['h0C7]=8'hC9;
    rom['h0C8]=8'hC0; rom['h0C9]=8'h2E; rom['h0CA]=8'h67; rom['h0CB]=8'h5D;
    rom['h0CC]=8'hD0; rom['h0CD]=8'h12; rom['h0CE]=8'hD0; rom['h0CF]=8'hC1;
    rom['h0D0]=8'hC0; rom['h0D1]=8'hFF; rom['h0D2]=8'hFF; rom['h0D3]=8'hFF;
    rom['h0D4]=8'hFF; rom['h0D5]=8'hFF; rom['h0D6]=8'hFF; rom['h0D7]=8'hFF;
    rom['h0D8]=8'hFF; rom['h0D9]=8'hFF; rom['h0DA]=8'hFF; rom['h0DB]=8'hFF;
    rom['h0DC]=8'hFF; rom['h0DD]=8'hFF; rom['h0DE]=8'hFF; rom['h0DF]=8'hFF;
    rom['h0E0]=8'hFF; rom['h0E1]=8'hFF; rom['h0E2]=8'hFF; rom['h0E3]=8'hFF;
    rom['h0E4]=8'hFF; rom['h0E5]=8'hFF; rom['h0E6]=8'hFF; rom['h0E7]=8'hFF;
    rom['h0E8]=8'hFF; rom['h0E9]=8'hFF; rom['h0EA]=8'hFF; rom['h0EB]=8'hFF;
    rom['h0EC]=8'hFF; rom['h0ED]=8'hFF; rom['h0EE]=8'hFF; rom['h0EF]=8'hFF;
    rom['h0F0]=8'hFF; rom['h0F1]=8'hFF; rom['h0F2]=8'hFF; rom['h0F3]=8'hFF;
    rom['h0F4]=8'hFF; rom['h0F5]=8'hFF; rom['h0F6]=8'hFF; rom['h0F7]=8'hFF;
    rom['h0F8]=8'hFF; rom['h0F9]=8'hFF; rom['h0FA]=8'hFF; rom['h0FB]=8'hFF;
    rom['h0FC]=8'hFF; rom['h0FD]=8'hFF; rom['h0FE]=8'hFF; rom['h0FF]=8'hFF;
    rom['h100]=8'h20; rom['h101]=8'h54; rom['h102]=8'h5E; rom['h103]=8'h00;
    rom['h104]=8'h22; rom['h105]=8'h00; rom['h106]=8'h20; rom['h107]=8'h78;
    rom['h108]=8'h56; rom['h109]=8'h5F; rom['h10A]=8'h20; rom['h10B]=8'h7A;
    rom['h10C]=8'h56; rom['h10D]=8'h5F; rom['h10E]=8'h20; rom['h10F]=8'h74;
    rom['h110]=8'h24; rom['h111]=8'h01; rom['h112]=8'h26; rom['h113]=8'h00;
    rom['h114]=8'h55; rom['h115]=8'hF9; rom['h116]=8'h20; rom['h117]=8'h78;
    rom['h118]=8'h56; rom['h119]=8'h6A; rom['h11A]=8'h5D; rom['h11B]=8'hF5;
    rom['h11C]=8'h14; rom['h11D]=8'h58; rom['h11E]=8'h20; rom['h11F]=8'h7C;
    rom['h120]=8'h5E; rom['h121]=8'h00; rom['h122]=8'h58; rom['h123]=8'hB0;
    rom['h124]=8'h20; rom['h125]=8'h7A; rom['h126]=8'h56; rom['h127]=8'h6A;
    rom['h128]=8'h58; rom['h129]=8'hB0; rom['h12A]=8'h5D; rom['h12B]=8'h53;
    rom['h12C]=8'h20; rom['h12D]=8'h83; rom['h12E]=8'h5E; rom['h12F]=8'h00;
    rom['h130]=8'h20; rom['h131]=8'h00; rom['h132]=8'h22; rom['h133]=8'h00;
    rom['h134]=8'h59; rom['h135]=8'hD9; rom['h136]=8'h55; rom['h137]=8'hDA;
    rom['h138]=8'h57; rom['h139]=8'hEC; rom['h13A]=8'h59; rom['h13B]=8'hFC;
    rom['h13C]=8'h5D; rom['h13D]=8'h5C; rom['h13E]=8'h22; rom['h13F]=8'h6C;
    rom['h140]=8'h55; rom['h141]=8'hB9; rom['h142]=8'h14; rom['h143]=8'h4E;
    rom['h144]=8'h20; rom['h145]=8'h8C; rom['h146]=8'h5E; rom['h147]=8'h00;
    rom['h148]=8'h22; rom['h149]=8'h6C; rom['h14A]=8'h58; rom['h14B]=8'h1D;
    rom['h14C]=8'h5D; rom['h14D]=8'h5C; rom['h14E]=8'h22; rom['h14F]=8'h00;
    rom['h150]=8'h20; rom['h151]=8'h78; rom['h152]=8'h56; rom['h153]=8'h5F;
    rom['h154]=8'h20; rom['h155]=8'h7A; rom['h156]=8'h56; rom['h157]=8'h5F;
    rom['h158]=8'h2E; rom['h159]=8'hFC; rom['h15A]=8'h2F; rom['h15B]=8'hEC;
    rom['h15C]=8'hB2; rom['h15D]=8'hED; rom['h15E]=8'hB3; rom['h15F]=8'h5D;
    rom['h160]=8'hF5; rom['h161]=8'h14; rom['h162]=8'h6F; rom['h163]=8'h20;
    rom['h164]=8'h88; rom['h165]=8'h5E; rom['h166]=8'h00; rom['h167]=8'hA2;
    rom['h168]=8'h5D; rom['h169]=8'h48; rom['h16A]=8'hA3; rom['h16B]=8'h5D;
    rom['h16C]=8'h48; rom['h16D]=8'h59; rom['h16E]=8'h39; rom['h16F]=8'h20;
    rom['h170]=8'h75; rom['h171]=8'h5E; rom['h172]=8'h00; rom['h173]=8'h20;
    rom['h174]=8'h6C; rom['h175]=8'h55; rom['h176]=8'h42; rom['h177]=8'h20;
    rom['h178]=8'h00; rom['h179]=8'h24; rom['h17A]=8'h00; rom['h17B]=8'h26;
    rom['h17C]=8'h00; rom['h17D]=8'h55; rom['h17E]=8'hF9; rom['h17F]=8'h5A;
    rom['h180]=8'h1D; rom['h181]=8'h59; rom['h182]=8'h06; rom['h183]=8'h2E;
    rom['h184]=8'h2E; rom['h185]=8'h5D; rom['h186]=8'hD0; rom['h187]=8'h1C;
    rom['h188]=8'h8B; rom['h189]=8'h40; rom['h18A]=8'h1B; rom['h18B]=8'h5D;
    rom['h18C]=8'h8C; rom['h18D]=8'h14; rom['h18E]=8'h91; rom['h18F]=8'h41;
    rom['h190]=8'hA5; rom['h191]=8'h20; rom['h192]=8'h6C; rom['h193]=8'h24;
    rom['h194]=8'h00; rom['h195]=8'h26; rom['h196]=8'h00; rom['h197]=8'h55;
    rom['h198]=8'hF9; rom['h199]=8'h20; rom['h19A]=8'h70; rom['h19B]=8'h24;
    rom['h19C]=8'h0D; rom['h19D]=8'h26; rom['h19E]=8'hFF; rom['h19F]=8'h55;
    rom['h1A0]=8'hF9; rom['h1A1]=8'h20; rom['h1A2]=8'h00; rom['h1A3]=8'h42;
    rom['h1A4]=8'h72; rom['h1A5]=8'h22; rom['h1A6]=8'hA0; rom['h1A7]=8'h5A;
    rom['h1A8]=8'h64; rom['h1A9]=8'h55; rom['h1AA]=8'hB9; rom['h1AB]=8'h1C;
    rom['h1AC]=8'hAF; rom['h1AD]=8'h42; rom['h1AE]=8'h14; rom['h1AF]=8'h55;
    rom['h1B0]=8'hCA; rom['h1B1]=8'h56; rom['h1B2]=8'h23; rom['h1B3]=8'h20;
    rom['h1B4]=8'h74; rom['h1B5]=8'hA6; rom['h1B6]=8'hB2; rom['h1B7]=8'hA7;
    rom['h1B8]=8'hB3; rom['h1B9]=8'h59; rom['h1BA]=8'h21; rom['h1BB]=8'h55;
    rom['h1BC]=8'hCA; rom['h1BD]=8'hA4; rom['h1BE]=8'hB2; rom['h1BF]=8'hA5;
    rom['h1C0]=8'hB3; rom['h1C1]=8'h59; rom['h1C2]=8'h21; rom['h1C3]=8'h55;
    rom['h1C4]=8'hCA; rom['h1C5]=8'hA0; rom['h1C6]=8'hB2; rom['h1C7]=8'hA1;
    rom['h1C8]=8'hB3; rom['h1C9]=8'h59; rom['h1CA]=8'hD9; rom['h1CB]=8'h55;
    rom['h1CC]=8'hCA; rom['h1CD]=8'h55; rom['h1CE]=8'hCA; rom['h1CF]=8'h20;
    rom['h1D0]=8'h00; rom['h1D1]=8'h59; rom['h1D2]=8'h06; rom['h1D3]=8'h5D;
    rom['h1D4]=8'hF5; rom['h1D5]=8'h14; rom['h1D6]=8'hE1; rom['h1D7]=8'h55;
    rom['h1D8]=8'hCA; rom['h1D9]=8'h20; rom['h1DA]=8'h74; rom['h1DB]=8'h59;
    rom['h1DC]=8'h21; rom['h1DD]=8'h55; rom['h1DE]=8'hCA; rom['h1DF]=8'h41;
    rom['h1E0]=8'hCF; rom['h1E1]=8'h20; rom['h1E2]=8'h74; rom['h1E3]=8'h22;
    rom['h1E4]=8'h00; rom['h1E5]=8'h59; rom['h1E6]=8'h21; rom['h1E7]=8'h55;
    rom['h1E8]=8'hCA; rom['h1E9]=8'h56; rom['h1EA]=8'h75; rom['h1EB]=8'h22;
    rom['h1EC]=8'hA0; rom['h1ED]=8'h59; rom['h1EE]=8'hFC; rom['h1EF]=8'hA2;
    rom['h1F0]=8'hB0; rom['h1F1]=8'hA3; rom['h1F2]=8'hB1; rom['h1F3]=8'hA6;
    rom['h1F4]=8'hB2; rom['h1F5]=8'hA7; rom['h1F6]=8'hB3; rom['h1F7]=8'h59;
    rom['h1F8]=8'h21; rom['h1F9]=8'h55; rom['h1FA]=8'hCA; rom['h1FB]=8'hA4;
    rom['h1FC]=8'hB2; rom['h1FD]=8'hA5; rom['h1FE]=8'hB3; rom['h1FF]=8'h59;
    rom['h200]=8'h21; rom['h201]=8'h41; rom['h202]=8'h73; rom['h203]=8'h59;
    rom['h204]=8'h06; rom['h205]=8'h55; rom['h206]=8'hCA; rom['h207]=8'hA2;
    rom['h208]=8'hB6; rom['h209]=8'hA3; rom['h20A]=8'hB7; rom['h20B]=8'h59;
    rom['h20C]=8'h06; rom['h20D]=8'h55; rom['h20E]=8'hCA; rom['h20F]=8'hA2;
    rom['h210]=8'hB4; rom['h211]=8'hA3; rom['h212]=8'hB5; rom['h213]=8'hC0;
    rom['h214]=8'h20; rom['h215]=8'h00; rom['h216]=8'h24; rom['h217]=8'h01;
    rom['h218]=8'h26; rom['h219]=8'h00; rom['h21A]=8'h55; rom['h21B]=8'hF9;
    rom['h21C]=8'h22; rom['h21D]=8'h74; rom['h21E]=8'h57; rom['h21F]=8'hC8;
    rom['h220]=8'h1A; rom['h221]=8'h24; rom['h222]=8'h41; rom['h223]=8'h16;
    rom['h224]=8'h52; rom['h225]=8'h03; rom['h226]=8'h22; rom['h227]=8'h6C;
    rom['h228]=8'h56; rom['h229]=8'h0E; rom['h22A]=8'h58; rom['h22B]=8'h1D;
    rom['h22C]=8'h5D; rom['h22D]=8'h53; rom['h22E]=8'h55; rom['h22F]=8'hCA;
    rom['h230]=8'h55; rom['h231]=8'hCA; rom['h232]=8'h57; rom['h233]=8'hEC;
    rom['h234]=8'h5D; rom['h235]=8'h5C; rom['h236]=8'h55; rom['h237]=8'hCA;
    rom['h238]=8'h42; rom['h239]=8'h1C; rom['h23A]=8'h20; rom['h23B]=8'h00;
    rom['h23C]=8'h24; rom['h23D]=8'h01; rom['h23E]=8'h26; rom['h23F]=8'h00;
    rom['h240]=8'h55; rom['h241]=8'hF9; rom['h242]=8'h52; rom['h243]=8'h03;
    rom['h244]=8'h20; rom['h245]=8'hA0; rom['h246]=8'h55; rom['h247]=8'hF9;
    rom['h248]=8'h22; rom['h249]=8'h6C; rom['h24A]=8'h57; rom['h24B]=8'hC8;
    rom['h24C]=8'h12; rom['h24D]=8'h5C; rom['h24E]=8'h20; rom['h24F]=8'h00;
    rom['h250]=8'h52; rom['h251]=8'h03; rom['h252]=8'h22; rom['h253]=8'h74;
    rom['h254]=8'h55; rom['h255]=8'hF9; rom['h256]=8'h57; rom['h257]=8'hC8;
    rom['h258]=8'h12; rom['h259]=8'h60; rom['h25A]=8'h42; rom['h25B]=8'h42;
    rom['h25C]=8'h55; rom['h25D]=8'h62; rom['h25E]=8'h42; rom['h25F]=8'h6A;
    rom['h260]=8'h41; rom['h261]=8'h16; rom['h262]=8'h20; rom['h263]=8'h00;
    rom['h264]=8'h52; rom['h265]=8'h03; rom['h266]=8'h20; rom['h267]=8'h6C;
    rom['h268]=8'h55; rom['h269]=8'hF9; rom['h26A]=8'h20; rom['h26B]=8'h00;
    rom['h26C]=8'h52; rom['h26D]=8'h03; rom['h26E]=8'h20; rom['h26F]=8'h70;
    rom['h270]=8'h55; rom['h271]=8'hF9; rom['h272]=8'h42; rom['h273]=8'h86;
    rom['h274]=8'h20; rom['h275]=8'h74; rom['h276]=8'h22; rom['h277]=8'h70;
    rom['h278]=8'h57; rom['h279]=8'hC8; rom['h27A]=8'h1A; rom['h27B]=8'h84;
    rom['h27C]=8'h14; rom['h27D]=8'h84; rom['h27E]=8'h20; rom['h27F]=8'h00;
    rom['h280]=8'h55; rom['h281]=8'h4F; rom['h282]=8'h42; rom['h283]=8'h62;
    rom['h284]=8'h41; rom['h285]=8'h16; rom['h286]=8'h20; rom['h287]=8'h00;
    rom['h288]=8'h55; rom['h289]=8'h1C; rom['h28A]=8'h59; rom['h28B]=8'h06;
    rom['h28C]=8'h5D; rom['h28D]=8'hF5; rom['h28E]=8'h1C; rom['h28F]=8'h92;
    rom['h290]=8'h42; rom['h291]=8'h74; rom['h292]=8'h55; rom['h293]=8'hCA;
    rom['h294]=8'h2E; rom['h295]=8'h3F; rom['h296]=8'h5D; rom['h297]=8'hD0;
    rom['h298]=8'h14; rom['h299]=8'h9C; rom['h29A]=8'h42; rom['h29B]=8'hBD;
    rom['h29C]=8'h59; rom['h29D]=8'h06; rom['h29E]=8'h2E; rom['h29F]=8'h24;
    rom['h2A0]=8'h5D; rom['h2A1]=8'hD0; rom['h2A2]=8'h1C; rom['h2A3]=8'hAB;
    rom['h2A4]=8'h55; rom['h2A5]=8'hCA; rom['h2A6]=8'hD1; rom['h2A7]=8'h53;
    rom['h2A8]=8'h39; rom['h2A9]=8'h43; rom['h2AA]=8'h44; rom['h2AB]=8'h2E;
    rom['h2AC]=8'h3F; rom['h2AD]=8'h5D; rom['h2AE]=8'hD0; rom['h2AF]=8'h1C;
    rom['h2B0]=8'hB8; rom['h2B1]=8'h55; rom['h2B2]=8'hCA; rom['h2B3]=8'hD2;
    rom['h2B4]=8'h53; rom['h2B5]=8'h39; rom['h2B6]=8'h43; rom['h2B7]=8'h44;
    rom['h2B8]=8'hD0; rom['h2B9]=8'h53; rom['h2BA]=8'h39; rom['h2BB]=8'h43;
    rom['h2BC]=8'h44; rom['h2BD]=8'h55; rom['h2BE]=8'hCA; rom['h2BF]=8'h59;
    rom['h2C0]=8'h5B; rom['h2C1]=8'h22; rom['h2C2]=8'h8C; rom['h2C3]=8'h24;
    rom['h2C4]=8'hDD; rom['h2C5]=8'h43; rom['h2C6]=8'h94; rom['h2C7]=8'h24;
    rom['h2C8]=8'h8C; rom['h2C9]=8'h59; rom['h2CA]=8'hA5; rom['h2CB]=8'h5D;
    rom['h2CC]=8'h9A; rom['h2CD]=8'h14; rom['h2CE]=8'hD5; rom['h2CF]=8'h55;
    rom['h2D0]=8'h2D; rom['h2D1]=8'h55; rom['h2D2]=8'h75; rom['h2D3]=8'h42;
    rom['h2D4]=8'h86; rom['h2D5]=8'h2E; rom['h2D6]=8'h3B; rom['h2D7]=8'h5D;
    rom['h2D8]=8'hD0; rom['h2D9]=8'h1C; rom['h2DA]=8'hE5; rom['h2DB]=8'h22;
    rom['h2DC]=8'h8C; rom['h2DD]=8'h55; rom['h2DE]=8'hB9; rom['h2DF]=8'h1C;
    rom['h2E0]=8'hE3; rom['h2E1]=8'h42; rom['h2E2]=8'h74; rom['h2E3]=8'h42;
    rom['h2E4]=8'h86; rom['h2E5]=8'h2E; rom['h2E6]=8'h23; rom['h2E7]=8'h5D;
    rom['h2E8]=8'hD0; rom['h2E9]=8'h1C; rom['h2EA]=8'hF9; rom['h2EB]=8'h22;
    rom['h2EC]=8'h8C; rom['h2ED]=8'h55; rom['h2EE]=8'hB9; rom['h2EF]=8'h14;
    rom['h2F0]=8'hF7; rom['h2F1]=8'h22; rom['h2F2]=8'h6C; rom['h2F3]=8'h55;
    rom['h2F4]=8'h75; rom['h2F5]=8'h42; rom['h2F6]=8'h3A; rom['h2F7]=8'h42;
    rom['h2F8]=8'h86; rom['h2F9]=8'h2E; rom['h2FA]=8'h21; rom['h2FB]=8'h5D;
    rom['h2FC]=8'hD0; rom['h2FD]=8'h00; rom['h2FE]=8'h00; rom['h2FF]=8'h00;
    rom['h300]=8'h00; rom['h301]=8'h14; rom['h302]=8'h05; rom['h303]=8'h43;
    rom['h304]=8'h11; rom['h305]=8'h20; rom['h306]=8'h94; rom['h307]=8'h22;
    rom['h308]=8'h6C; rom['h309]=8'h55; rom['h30A]=8'h4F; rom['h30B]=8'h55;
    rom['h30C]=8'hCA; rom['h30D]=8'h20; rom['h30E]=8'h00; rom['h30F]=8'h42;
    rom['h310]=8'hEB; rom['h311]=8'h2E; rom['h312]=8'h26; rom['h313]=8'h5D;
    rom['h314]=8'hD0; rom['h315]=8'h1C; rom['h316]=8'h1D; rom['h317]=8'h22;
    rom['h318]=8'h74; rom['h319]=8'h55; rom['h31A]=8'h75; rom['h31B]=8'h42;
    rom['h31C]=8'h86; rom['h31D]=8'h2E; rom['h31E]=8'h24; rom['h31F]=8'h5D;
    rom['h320]=8'hD0; rom['h321]=8'h1C; rom['h322]=8'h2D; rom['h323]=8'hA4;
    rom['h324]=8'hB0; rom['h325]=8'hA5; rom['h326]=8'hB1; rom['h327]=8'h56;
    rom['h328]=8'h6A; rom['h329]=8'h5D; rom['h32A]=8'h28; rom['h32B]=8'h42;
    rom['h32C]=8'h86; rom['h32D]=8'h20; rom['h32E]=8'h7A; rom['h32F]=8'h56;
    rom['h330]=8'h5F; rom['h331]=8'h20; rom['h332]=8'h78; rom['h333]=8'h22;
    rom['h334]=8'hE0; rom['h335]=8'h56; rom['h336]=8'h5F; rom['h337]=8'h41;
    rom['h338]=8'h16; rom['h339]=8'h2E; rom['h33A]=8'h7E; rom['h33B]=8'h2F;
    rom['h33C]=8'hE0; rom['h33D]=8'hC0; rom['h33E]=8'h2E; rom['h33F]=8'h7E;
    rom['h340]=8'h2F; rom['h341]=8'hE9; rom['h342]=8'hB5; rom['h343]=8'hC0;
    rom['h344]=8'h55; rom['h345]=8'hCA; rom['h346]=8'h59; rom['h347]=8'h06;
    rom['h348]=8'h5D; rom['h349]=8'hF5; rom['h34A]=8'h1C; rom['h34B]=8'h4E;
    rom['h34C]=8'h43; rom['h34D]=8'h8C; rom['h34E]=8'h2E; rom['h34F]=8'h22;
    rom['h350]=8'h5D; rom['h351]=8'hD0; rom['h352]=8'h1C; rom['h353]=8'h56;
    rom['h354]=8'h43; rom['h355]=8'h78; rom['h356]=8'h22; rom['h357]=8'h8C;
    rom['h358]=8'h24; rom['h359]=8'hE7; rom['h35A]=8'h43; rom['h35B]=8'h94;
    rom['h35C]=8'h53; rom['h35D]=8'h3E; rom['h35E]=8'hF0; rom['h35F]=8'hD1;
    rom['h360]=8'h95; rom['h361]=8'h1C; rom['h362]=8'h6B; rom['h363]=8'h20;
    rom['h364]=8'h8C; rom['h365]=8'h56; rom['h366]=8'h6A; rom['h367]=8'h58;
    rom['h368]=8'hB0; rom['h369]=8'h43; rom['h36A]=8'h92; rom['h36B]=8'hF0;
    rom['h36C]=8'hD2; rom['h36D]=8'h95; rom['h36E]=8'h1C; rom['h36F]=8'h74;
    rom['h370]=8'h58; rom['h371]=8'h8D; rom['h372]=8'h43; rom['h373]=8'h92;
    rom['h374]=8'h58; rom['h375]=8'h1D; rom['h376]=8'h43; rom['h377]=8'h92;
    rom['h378]=8'h55; rom['h379]=8'hCA; rom['h37A]=8'h57; rom['h37B]=8'hF4;
    rom['h37C]=8'h59; rom['h37D]=8'h06; rom['h37E]=8'h2E; rom['h37F]=8'h3B;
    rom['h380]=8'h5D; rom['h381]=8'hD0; rom['h382]=8'h14; rom['h383]=8'h88;
    rom['h384]=8'h5D; rom['h385]=8'h5C; rom['h386]=8'h43; rom['h387]=8'h92;
    rom['h388]=8'h55; rom['h389]=8'hCA; rom['h38A]=8'h43; rom['h38B]=8'h92;
    rom['h38C]=8'h20; rom['h38D]=8'h78; rom['h38E]=8'h22; rom['h38F]=8'hA0;
    rom['h390]=8'h41; rom['h391]=8'h16; rom['h392]=8'h42; rom['h393]=8'h86;
    rom['h394]=8'h59; rom['h395]=8'h73; rom['h396]=8'h59; rom['h397]=8'h5B;
    rom['h398]=8'h20; rom['h399]=8'h00; rom['h39A]=8'h59; rom['h39B]=8'h06;
    rom['h39C]=8'h5D; rom['h39D]=8'hF5; rom['h39E]=8'h1C; rom['h39F]=8'hA8;
    rom['h3A0]=8'h20; rom['h3A1]=8'h78; rom['h3A2]=8'h22; rom['h3A3]=8'hE1;
    rom['h3A4]=8'h56; rom['h3A5]=8'h5F; rom['h3A6]=8'h41; rom['h3A7]=8'h16;
    rom['h3A8]=8'h22; rom['h3A9]=8'h80; rom['h3AA]=8'h24; rom['h3AB]=8'hDF;
    rom['h3AC]=8'h44; rom['h3AD]=8'h50; rom['h3AE]=8'h20; rom['h3AF]=8'h00;
    rom['h3B0]=8'h22; rom['h3B1]=8'h80; rom['h3B2]=8'h59; rom['h3B3]=8'hD9;
    rom['h3B4]=8'h59; rom['h3B5]=8'h06; rom['h3B6]=8'h5D; rom['h3B7]=8'hF5;
    rom['h3B8]=8'h1C; rom['h3B9]=8'hBC; rom['h3BA]=8'h44; rom['h3BB]=8'h40;
    rom['h3BC]=8'h55; rom['h3BD]=8'hCA; rom['h3BE]=8'h2E; rom['h3BF]=8'h29;
    rom['h3C0]=8'h5D; rom['h3C1]=8'hD0; rom['h3C2]=8'h1C; rom['h3C3]=8'hC6;
    rom['h3C4]=8'h44; rom['h3C5]=8'h40; rom['h3C6]=8'h2E; rom['h3C7]=8'h20;
    rom['h3C8]=8'h5D; rom['h3C9]=8'hD0; rom['h3CA]=8'h1C; rom['h3CB]=8'hCE;
    rom['h3CC]=8'h44; rom['h3CD]=8'h40; rom['h3CE]=8'h59; rom['h3CF]=8'h5B;
    rom['h3D0]=8'h22; rom['h3D1]=8'h84; rom['h3D2]=8'h24; rom['h3D3]=8'hE1;
    rom['h3D4]=8'h44; rom['h3D5]=8'h50; rom['h3D6]=8'h59; rom['h3D7]=8'hBF;
    rom['h3D8]=8'h22; rom['h3D9]=8'h80; rom['h3DA]=8'h59; rom['h3DB]=8'hFC;
    rom['h3DC]=8'h20; rom['h3DD]=8'h80; rom['h3DE]=8'h22; rom['h3DF]=8'h84;
    rom['h3E0]=8'h2E; rom['h3E1]=8'h2B; rom['h3E2]=8'h5D; rom['h3E3]=8'hE9;
    rom['h3E4]=8'h1C; rom['h3E5]=8'hEA; rom['h3E6]=8'h56; rom['h3E7]=8'hC0;
    rom['h3E8]=8'h43; rom['h3E9]=8'hAE; rom['h3EA]=8'h2E; rom['h3EB]=8'h2D;
    rom['h3EC]=8'h5D; rom['h3ED]=8'hE9; rom['h3EE]=8'h1C; rom['h3EF]=8'hF4;
    rom['h3F0]=8'h56; rom['h3F1]=8'hD5; rom['h3F2]=8'h43; rom['h3F3]=8'hAE;
    rom['h3F4]=8'h2E; rom['h3F5]=8'h2A; rom['h3F6]=8'h5D; rom['h3F7]=8'hE9;
    rom['h3F8]=8'h1C; rom['h3F9]=8'hFE; rom['h3FA]=8'h56; rom['h3FB]=8'hFE;
    rom['h3FC]=8'h43; rom['h3FD]=8'hAE; rom['h3FE]=8'h2E; rom['h3FF]=8'h2F;
    rom['h400]=8'h5D; rom['h401]=8'hE9; rom['h402]=8'h00; rom['h403]=8'h00;
    rom['h404]=8'h1C; rom['h405]=8'h0A; rom['h406]=8'h57; rom['h407]=8'h21;
    rom['h408]=8'h43; rom['h409]=8'hAE; rom['h40A]=8'h2E; rom['h40B]=8'h3D;
    rom['h40C]=8'h5D; rom['h40D]=8'hE9; rom['h40E]=8'h1C; rom['h40F]=8'h1E;
    rom['h410]=8'h57; rom['h411]=8'hC8; rom['h412]=8'h14; rom['h413]=8'h18;
    rom['h414]=8'h55; rom['h415]=8'h42; rom['h416]=8'h43; rom['h417]=8'hAE;
    rom['h418]=8'h22; rom['h419]=8'h01; rom['h41A]=8'h56; rom['h41B]=8'h38;
    rom['h41C]=8'h43; rom['h41D]=8'hAE; rom['h41E]=8'h2E; rom['h41F]=8'h3C;
    rom['h420]=8'h5D; rom['h421]=8'hE9; rom['h422]=8'h1C; rom['h423]=8'h2A;
    rom['h424]=8'h57; rom['h425]=8'hC8; rom['h426]=8'h1A; rom['h427]=8'h18;
    rom['h428]=8'h44; rom['h429]=8'h14; rom['h42A]=8'h2E; rom['h42B]=8'h3E;
    rom['h42C]=8'h5D; rom['h42D]=8'hE9; rom['h42E]=8'h1C; rom['h42F]=8'h36;
    rom['h430]=8'h57; rom['h431]=8'hC8; rom['h432]=8'h1A; rom['h433]=8'h14;
    rom['h434]=8'h44; rom['h435]=8'h18; rom['h436]=8'h20; rom['h437]=8'h78;
    rom['h438]=8'h22; rom['h439]=8'hE2; rom['h43A]=8'h22; rom['h43B]=8'h80;
    rom['h43C]=8'h59; rom['h43D]=8'hD9; rom['h43E]=8'h41; rom['h43F]=8'h16;
    rom['h440]=8'h22; rom['h441]=8'hA0; rom['h442]=8'h59; rom['h443]=8'hFC;
    rom['h444]=8'h59; rom['h445]=8'hA5; rom['h446]=8'h20; rom['h447]=8'hA0;
    rom['h448]=8'h55; rom['h449]=8'h62; rom['h44A]=8'h20; rom['h44B]=8'h00;
    rom['h44C]=8'h59; rom['h44D]=8'hBF; rom['h44E]=8'h4B; rom['h44F]=8'hD0;
    rom['h450]=8'h59; rom['h451]=8'h73; rom['h452]=8'h59; rom['h453]=8'h5B;
    rom['h454]=8'h20; rom['h455]=8'h00; rom['h456]=8'h59; rom['h457]=8'h06;
    rom['h458]=8'h2E; rom['h459]=8'h28; rom['h45A]=8'h5D; rom['h45B]=8'hD0;
    rom['h45C]=8'h1C; rom['h45D]=8'h68; rom['h45E]=8'h55; rom['h45F]=8'hCA;
    rom['h460]=8'h24; rom['h461]=8'hE3; rom['h462]=8'h22; rom['h463]=8'h88;
    rom['h464]=8'h43; rom['h465]=8'h94; rom['h466]=8'h45; rom['h467]=8'h10;
    rom['h468]=8'h24; rom['h469]=8'h88; rom['h46A]=8'h2E; rom['h46B]=8'h2D;
    rom['h46C]=8'h5D; rom['h46D]=8'hD0; rom['h46E]=8'h1C; rom['h46F]=8'h80;
    rom['h470]=8'h55; rom['h471]=8'hCA; rom['h472]=8'h24; rom['h473]=8'hE5;
    rom['h474]=8'h22; rom['h475]=8'h88; rom['h476]=8'h44; rom['h477]=8'h50;
    rom['h478]=8'h20; rom['h479]=8'h88; rom['h47A]=8'h55; rom['h47B]=8'hEB;
    rom['h47C]=8'h55; rom['h47D]=8'hCA; rom['h47E]=8'h45; rom['h47F]=8'h10;
    rom['h480]=8'h5D; rom['h481]=8'h8C; rom['h482]=8'h14; rom['h483]=8'h8A;
    rom['h484]=8'h22; rom['h485]=8'h88; rom['h486]=8'h5A; rom['h487]=8'h64;
    rom['h488]=8'h45; rom['h489]=8'h10; rom['h48A]=8'h5D; rom['h48B]=8'h9A;
    rom['h48C]=8'h14; rom['h48D]=8'h94; rom['h48E]=8'h55; rom['h48F]=8'h2D;
    rom['h490]=8'h55; rom['h491]=8'h9B; rom['h492]=8'h45; rom['h493]=8'h0E;
    rom['h494]=8'h2E; rom['h495]=8'h25; rom['h496]=8'h5D; rom['h497]=8'hD0;
    rom['h498]=8'h1C; rom['h499]=8'hA0; rom['h49A]=8'h22; rom['h49B]=8'h90;
    rom['h49C]=8'h55; rom['h49D]=8'h9B; rom['h49E]=8'h45; rom['h49F]=8'h0E;
    rom['h4A0]=8'h2E; rom['h4A1]=8'h23; rom['h4A2]=8'h5D; rom['h4A3]=8'hD0;
    rom['h4A4]=8'h1C; rom['h4A5]=8'hAC; rom['h4A6]=8'h22; rom['h4A7]=8'h6C;
    rom['h4A8]=8'h55; rom['h4A9]=8'h9B; rom['h4AA]=8'h45; rom['h4AB]=8'h0E;
    rom['h4AC]=8'h2E; rom['h4AD]=8'h21; rom['h4AE]=8'h5D; rom['h4AF]=8'hD0;
    rom['h4B0]=8'h1C; rom['h4B1]=8'hB8; rom['h4B2]=8'h22; rom['h4B3]=8'h94;
    rom['h4B4]=8'h55; rom['h4B5]=8'h9B; rom['h4B6]=8'h45; rom['h4B7]=8'h0E;
    rom['h4B8]=8'h2E; rom['h4B9]=8'h27; rom['h4BA]=8'h5D; rom['h4BB]=8'hD0;
    rom['h4BC]=8'h1C; rom['h4BD]=8'hC4; rom['h4BE]=8'h22; rom['h4BF]=8'h98;
    rom['h4C0]=8'h55; rom['h4C1]=8'h9B; rom['h4C2]=8'h45; rom['h4C3]=8'h0E;
    rom['h4C4]=8'h2E; rom['h4C5]=8'h26; rom['h4C6]=8'h5D; rom['h4C7]=8'hD0;
    rom['h4C8]=8'h1C; rom['h4C9]=8'hD0; rom['h4CA]=8'h22; rom['h4CB]=8'h74;
    rom['h4CC]=8'h55; rom['h4CD]=8'h9B; rom['h4CE]=8'h45; rom['h4CF]=8'h0E;
    rom['h4D0]=8'h2E; rom['h4D1]=8'h24; rom['h4D2]=8'h5D; rom['h4D3]=8'hD0;
    rom['h4D4]=8'h1C; rom['h4D5]=8'hE0; rom['h4D6]=8'h5D; rom['h4D7]=8'h00;
    rom['h4D8]=8'h20; rom['h4D9]=8'h88; rom['h4DA]=8'h56; rom['h4DB]=8'h38;
    rom['h4DC]=8'h20; rom['h4DD]=8'h00; rom['h4DE]=8'h45; rom['h4DF]=8'h0E;
    rom['h4E0]=8'h2E; rom['h4E1]=8'h3F; rom['h4E2]=8'h5D; rom['h4E3]=8'hD0;
    rom['h4E4]=8'h14; rom['h4E5]=8'hE8; rom['h4E6]=8'h45; rom['h4E7]=8'h02;
    rom['h4E8]=8'h20; rom['h4E9]=8'h00; rom['h4EA]=8'h22; rom['h4EB]=8'h00;
    rom['h4EC]=8'h59; rom['h4ED]=8'hD9; rom['h4EE]=8'h24; rom['h4EF]=8'h00;
    rom['h4F0]=8'h26; rom['h4F1]=8'h00; rom['h4F2]=8'h55; rom['h4F3]=8'hF9;
    rom['h4F4]=8'h5A; rom['h4F5]=8'h1D; rom['h4F6]=8'h22; rom['h4F7]=8'h88;
    rom['h4F8]=8'h24; rom['h4F9]=8'hE9; rom['h4FA]=8'h43; rom['h4FB]=8'h94;
    rom['h4FC]=8'h22; rom['h4FD]=8'h00; rom['h4FE]=8'h59; rom['h4FF]=8'hFC;
    rom['h500]=8'h45; rom['h501]=8'h0E; rom['h502]=8'h20; rom['h503]=8'h7A;
    rom['h504]=8'h56; rom['h505]=8'h5F; rom['h506]=8'h22; rom['h507]=8'hF0;
    rom['h508]=8'h20; rom['h509]=8'h78; rom['h50A]=8'h56; rom['h50B]=8'h5F;
    rom['h50C]=8'h41; rom['h50D]=8'h16; rom['h50E]=8'h55; rom['h50F]=8'hCA;
    rom['h510]=8'h59; rom['h511]=8'hA5; rom['h512]=8'h20; rom['h513]=8'h88;
    rom['h514]=8'h55; rom['h515]=8'h62; rom['h516]=8'h20; rom['h517]=8'h00;
    rom['h518]=8'h59; rom['h519]=8'hBF; rom['h51A]=8'h4B; rom['h51B]=8'hD0;
    rom['h51C]=8'h59; rom['h51D]=8'h5B; rom['h51E]=8'h59; rom['h51F]=8'h06;
    rom['h520]=8'h2E; rom['h521]=8'h20; rom['h522]=8'h5D; rom['h523]=8'hD0;
    rom['h524]=8'h1C; rom['h525]=8'h2A; rom['h526]=8'h55; rom['h527]=8'hCA;
    rom['h528]=8'h45; rom['h529]=8'h1E; rom['h52A]=8'h59; rom['h52B]=8'hA5;
    rom['h52C]=8'hC0; rom['h52D]=8'hF0; rom['h52E]=8'hA2; rom['h52F]=8'hF6;
    rom['h530]=8'hF7; rom['h531]=8'hF5; rom['h532]=8'hF5; rom['h533]=8'hB2;
    rom['h534]=8'hA3; rom['h535]=8'hF6; rom['h536]=8'hF1; rom['h537]=8'hF6;
    rom['h538]=8'hF1; rom['h539]=8'h82; rom['h53A]=8'hB2; rom['h53B]=8'hF0;
    rom['h53C]=8'hA3; rom['h53D]=8'hF5; rom['h53E]=8'hF1; rom['h53F]=8'hF5;
    rom['h540]=8'hB3; rom['h541]=8'hC0; rom['h542]=8'hA1; rom['h543]=8'hBF;
    rom['h544]=8'hDC; rom['h545]=8'hBE; rom['h546]=8'hF0; rom['h547]=8'h21;
    rom['h548]=8'hE0; rom['h549]=8'h61; rom['h54A]=8'h7E; rom['h54B]=8'h47;
    rom['h54C]=8'hAF; rom['h54D]=8'hB1; rom['h54E]=8'hC0; rom['h54F]=8'hA1;
    rom['h550]=8'hBF; rom['h551]=8'hA3; rom['h552]=8'hBD; rom['h553]=8'hDC;
    rom['h554]=8'hBE; rom['h555]=8'h23; rom['h556]=8'hE9; rom['h557]=8'h21;
    rom['h558]=8'hE0; rom['h559]=8'h61; rom['h55A]=8'h63; rom['h55B]=8'h7E;
    rom['h55C]=8'h55; rom['h55D]=8'hAF; rom['h55E]=8'hB1; rom['h55F]=8'hAD;
    rom['h560]=8'hB3; rom['h561]=8'hC0; rom['h562]=8'hA1; rom['h563]=8'hBF;
    rom['h564]=8'hA3; rom['h565]=8'hBD; rom['h566]=8'hDC; rom['h567]=8'hBE;
    rom['h568]=8'h21; rom['h569]=8'hE9; rom['h56A]=8'h23; rom['h56B]=8'hE0;
    rom['h56C]=8'h61; rom['h56D]=8'h63; rom['h56E]=8'h7E; rom['h56F]=8'h68;
    rom['h570]=8'hAF; rom['h571]=8'hB1; rom['h572]=8'hAD; rom['h573]=8'hB3;
    rom['h574]=8'hC0; rom['h575]=8'hA5; rom['h576]=8'hBF; rom['h577]=8'hA3;
    rom['h578]=8'hBD; rom['h579]=8'hDC; rom['h57A]=8'hBE; rom['h57B]=8'h25;
    rom['h57C]=8'hE9; rom['h57D]=8'h23; rom['h57E]=8'hE0; rom['h57F]=8'h65;
    rom['h580]=8'h63; rom['h581]=8'h7E; rom['h582]=8'h7B; rom['h583]=8'hAF;
    rom['h584]=8'hB5; rom['h585]=8'hAD; rom['h586]=8'hB3; rom['h587]=8'hC0;
    rom['h588]=8'hA1; rom['h589]=8'hBF; rom['h58A]=8'hA5; rom['h58B]=8'hBD;
    rom['h58C]=8'hDC; rom['h58D]=8'hBE; rom['h58E]=8'h21; rom['h58F]=8'hE9;
    rom['h590]=8'h25; rom['h591]=8'hE0; rom['h592]=8'h61; rom['h593]=8'h65;
    rom['h594]=8'h7E; rom['h595]=8'h8E; rom['h596]=8'hAF; rom['h597]=8'hB1;
    rom['h598]=8'hAD; rom['h599]=8'hB5; rom['h59A]=8'hC0; rom['h59B]=8'hA3;
    rom['h59C]=8'hBF; rom['h59D]=8'hA5; rom['h59E]=8'hBD; rom['h59F]=8'hDC;
    rom['h5A0]=8'hBE; rom['h5A1]=8'h23; rom['h5A2]=8'hE9; rom['h5A3]=8'h25;
    rom['h5A4]=8'hE0; rom['h5A5]=8'h63; rom['h5A6]=8'h65; rom['h5A7]=8'h7E;
    rom['h5A8]=8'hA1; rom['h5A9]=8'hAF; rom['h5AA]=8'hB3; rom['h5AB]=8'hAD;
    rom['h5AC]=8'hB5; rom['h5AD]=8'hC0; rom['h5AE]=8'hA1; rom['h5AF]=8'hBF;
    rom['h5B0]=8'h61; rom['h5B1]=8'h61; rom['h5B2]=8'h61; rom['h5B3]=8'h21;
    rom['h5B4]=8'hE9; rom['h5B5]=8'hF5; rom['h5B6]=8'hAF; rom['h5B7]=8'hB1;
    rom['h5B8]=8'hC0; rom['h5B9]=8'hA3; rom['h5BA]=8'hBF; rom['h5BB]=8'hDC;
    rom['h5BC]=8'hBE; rom['h5BD]=8'h23; rom['h5BE]=8'hE9; rom['h5BF]=8'h1C;
    rom['h5C0]=8'hC7; rom['h5C1]=8'h63; rom['h5C2]=8'h7E; rom['h5C3]=8'hBD;
    rom['h5C4]=8'hAF; rom['h5C5]=8'hB3; rom['h5C6]=8'hC0; rom['h5C7]=8'hAF;
    rom['h5C8]=8'hB3; rom['h5C9]=8'hC1; rom['h5CA]=8'hA1; rom['h5CB]=8'hBF;
    rom['h5CC]=8'hDC; rom['h5CD]=8'hBE; rom['h5CE]=8'h21; rom['h5CF]=8'hE9;
    rom['h5D0]=8'hF2; rom['h5D1]=8'hE0; rom['h5D2]=8'h1C; rom['h5D3]=8'hD7;
    rom['h5D4]=8'h61; rom['h5D5]=8'h7E; rom['h5D6]=8'hCE; rom['h5D7]=8'hAF;
    rom['h5D8]=8'hB1; rom['h5D9]=8'hC0; rom['h5DA]=8'hA1; rom['h5DB]=8'hBF;
    rom['h5DC]=8'hDC; rom['h5DD]=8'hBE; rom['h5DE]=8'hF1; rom['h5DF]=8'h21;
    rom['h5E0]=8'hE9; rom['h5E1]=8'hF8; rom['h5E2]=8'hE0; rom['h5E3]=8'h12;
    rom['h5E4]=8'hE8; rom['h5E5]=8'h61; rom['h5E6]=8'h7E; rom['h5E7]=8'hDF;
    rom['h5E8]=8'hAF; rom['h5E9]=8'hB1; rom['h5EA]=8'hC0; rom['h5EB]=8'hA1;
    rom['h5EC]=8'hBF; rom['h5ED]=8'hDC; rom['h5EE]=8'hBE; rom['h5EF]=8'h21;
    rom['h5F0]=8'hE9; rom['h5F1]=8'hF4; rom['h5F2]=8'hE0; rom['h5F3]=8'h61;
    rom['h5F4]=8'h7E; rom['h5F5]=8'hEF; rom['h5F6]=8'hAF; rom['h5F7]=8'hB1;
    rom['h5F8]=8'hC0; rom['h5F9]=8'h21; rom['h5FA]=8'hA7; rom['h5FB]=8'hE0;
    rom['h5FC]=8'h61; rom['h5FD]=8'h21; rom['h5FE]=8'hA6; rom['h5FF]=8'hE0;
    rom['h600]=8'h61; rom['h601]=8'h21; rom['h602]=8'hA5; rom['h603]=8'hE0;
    rom['h604]=8'h61; rom['h605]=8'h21; rom['h606]=8'hA4; rom['h607]=8'hE0;
    rom['h608]=8'hA1; rom['h609]=8'hF8; rom['h60A]=8'hF8; rom['h60B]=8'hF8;
    rom['h60C]=8'hB1; rom['h60D]=8'hC0; rom['h60E]=8'h23; rom['h60F]=8'hA7;
    rom['h610]=8'hE0; rom['h611]=8'h63; rom['h612]=8'h23; rom['h613]=8'hA6;
    rom['h614]=8'hE0; rom['h615]=8'h63; rom['h616]=8'h23; rom['h617]=8'hA5;
    rom['h618]=8'hE0; rom['h619]=8'h63; rom['h61A]=8'h23; rom['h61B]=8'hA4;
    rom['h61C]=8'hE0; rom['h61D]=8'hA3; rom['h61E]=8'hF8; rom['h61F]=8'hF8;
    rom['h620]=8'hF8; rom['h621]=8'hB3; rom['h622]=8'hC0; rom['h623]=8'h23;
    rom['h624]=8'hE9; rom['h625]=8'hB7; rom['h626]=8'h63; rom['h627]=8'h23;
    rom['h628]=8'hE9; rom['h629]=8'hB6; rom['h62A]=8'h63; rom['h62B]=8'h23;
    rom['h62C]=8'hE9; rom['h62D]=8'hB5; rom['h62E]=8'h63; rom['h62F]=8'h23;
    rom['h630]=8'hE9; rom['h631]=8'hB4; rom['h632]=8'hA3; rom['h633]=8'hF8;
    rom['h634]=8'hF8; rom['h635]=8'hF8; rom['h636]=8'hB3; rom['h637]=8'hC0;
    rom['h638]=8'h21; rom['h639]=8'hA3; rom['h63A]=8'hE0; rom['h63B]=8'h61;
    rom['h63C]=8'h21; rom['h63D]=8'hA2; rom['h63E]=8'hE0; rom['h63F]=8'hF0;
    rom['h640]=8'h61; rom['h641]=8'h21; rom['h642]=8'hE0; rom['h643]=8'h61;
    rom['h644]=8'h21; rom['h645]=8'hE0; rom['h646]=8'hA1; rom['h647]=8'hF8;
    rom['h648]=8'hF8; rom['h649]=8'hF8; rom['h64A]=8'hB1; rom['h64B]=8'hC0;
    rom['h64C]=8'h2E; rom['h64D]=8'h7D; rom['h64E]=8'h2F; rom['h64F]=8'hF0;
    rom['h650]=8'hE0; rom['h651]=8'hC0; rom['h652]=8'h2E; rom['h653]=8'h7D;
    rom['h654]=8'h2F; rom['h655]=8'hE9; rom['h656]=8'hF4; rom['h657]=8'hE0;
    rom['h658]=8'hC0; rom['h659]=8'h2E; rom['h65A]=8'h7D; rom['h65B]=8'h2F;
    rom['h65C]=8'hE9; rom['h65D]=8'hF6; rom['h65E]=8'hC0; rom['h65F]=8'h21;
    rom['h660]=8'hA3; rom['h661]=8'hE0; rom['h662]=8'h61; rom['h663]=8'h21;
    rom['h664]=8'hA2; rom['h665]=8'hE0; rom['h666]=8'hA1; rom['h667]=8'hF8;
    rom['h668]=8'hB1; rom['h669]=8'hC0; rom['h66A]=8'h21; rom['h66B]=8'hE9;
    rom['h66C]=8'hB3; rom['h66D]=8'h61; rom['h66E]=8'h21; rom['h66F]=8'hE9;
    rom['h670]=8'hB2; rom['h671]=8'hA1; rom['h672]=8'hF8; rom['h673]=8'hB1;
    rom['h674]=8'hC0; rom['h675]=8'h21; rom['h676]=8'hE9; rom['h677]=8'hB7;
    rom['h678]=8'h61; rom['h679]=8'h21; rom['h67A]=8'hE9; rom['h67B]=8'hB6;
    rom['h67C]=8'h61; rom['h67D]=8'h21; rom['h67E]=8'hE9; rom['h67F]=8'hB5;
    rom['h680]=8'h61; rom['h681]=8'h21; rom['h682]=8'hE9; rom['h683]=8'hB4;
    rom['h684]=8'hA1; rom['h685]=8'hF8; rom['h686]=8'hF8; rom['h687]=8'hF8;
    rom['h688]=8'hB1; rom['h689]=8'hC0; rom['h68A]=8'hA1; rom['h68B]=8'hBF;
    rom['h68C]=8'hDC; rom['h68D]=8'hBE; rom['h68E]=8'hF1; rom['h68F]=8'h21;
    rom['h690]=8'hE9; rom['h691]=8'hF5; rom['h692]=8'hE0; rom['h693]=8'h61;
    rom['h694]=8'h7E; rom['h695]=8'h8F; rom['h696]=8'hAF; rom['h697]=8'hB1;
    rom['h698]=8'hC0; rom['h699]=8'hA3; rom['h69A]=8'hBF; rom['h69B]=8'hDC;
    rom['h69C]=8'hBE; rom['h69D]=8'hF1; rom['h69E]=8'h23; rom['h69F]=8'hE9;
    rom['h6A0]=8'hF5; rom['h6A1]=8'hE0; rom['h6A2]=8'h63; rom['h6A3]=8'h7E;
    rom['h6A4]=8'h9E; rom['h6A5]=8'hAF; rom['h6A6]=8'hB3; rom['h6A7]=8'hC0;
    rom['h6A8]=8'h65; rom['h6A9]=8'h65; rom['h6AA]=8'h65; rom['h6AB]=8'hDC;
    rom['h6AC]=8'hBE; rom['h6AD]=8'hF0; rom['h6AE]=8'hBF; rom['h6AF]=8'hAF;
    rom['h6B0]=8'hF6; rom['h6B1]=8'h25; rom['h6B2]=8'hE9; rom['h6B3]=8'hF6;
    rom['h6B4]=8'hE0; rom['h6B5]=8'hF7; rom['h6B6]=8'hBF; rom['h6B7]=8'hA5;
    rom['h6B8]=8'hF8; rom['h6B9]=8'hB5; rom['h6BA]=8'h7E; rom['h6BB]=8'hAF;
    rom['h6BC]=8'h65; rom['h6BD]=8'hAF; rom['h6BE]=8'hF6; rom['h6BF]=8'hC0;
    rom['h6C0]=8'hA1; rom['h6C1]=8'hBF; rom['h6C2]=8'hA3; rom['h6C3]=8'hBD;
    rom['h6C4]=8'hDC; rom['h6C5]=8'hBE; rom['h6C6]=8'hF1; rom['h6C7]=8'h23;
    rom['h6C8]=8'hE9; rom['h6C9]=8'h21; rom['h6CA]=8'hEB; rom['h6CB]=8'hE0;
    rom['h6CC]=8'h61; rom['h6CD]=8'h63; rom['h6CE]=8'h7E; rom['h6CF]=8'hC7;
    rom['h6D0]=8'hAF; rom['h6D1]=8'hB1; rom['h6D2]=8'hAD; rom['h6D3]=8'hB3;
    rom['h6D4]=8'hC0; rom['h6D5]=8'hA1; rom['h6D6]=8'hBF; rom['h6D7]=8'hA3;
    rom['h6D8]=8'hBD; rom['h6D9]=8'hDC; rom['h6DA]=8'hBE; rom['h6DB]=8'hFA;
    rom['h6DC]=8'hF3; rom['h6DD]=8'h21; rom['h6DE]=8'hE9; rom['h6DF]=8'h23;
    rom['h6E0]=8'hE8; rom['h6E1]=8'h21; rom['h6E2]=8'hE0; rom['h6E3]=8'h61;
    rom['h6E4]=8'h63; rom['h6E5]=8'h7E; rom['h6E6]=8'hDC; rom['h6E7]=8'hAF;
    rom['h6E8]=8'hB1; rom['h6E9]=8'hAD; rom['h6EA]=8'hB3; rom['h6EB]=8'hC0;
    rom['h6EC]=8'hA6; rom['h6ED]=8'hB7; rom['h6EE]=8'hA5; rom['h6EF]=8'hB6;
    rom['h6F0]=8'hA4; rom['h6F1]=8'hB5; rom['h6F2]=8'hF0; rom['h6F3]=8'hB4;
    rom['h6F4]=8'hC0; rom['h6F5]=8'hA5; rom['h6F6]=8'hB4; rom['h6F7]=8'hA6;
    rom['h6F8]=8'hB5; rom['h6F9]=8'hA7; rom['h6FA]=8'hB6; rom['h6FB]=8'hF0;
    rom['h6FC]=8'hB7; rom['h6FD]=8'hC0; rom['h6FE]=8'h59; rom['h6FF]=8'h5B;
    rom['h700]=8'h59; rom['h701]=8'h73; rom['h702]=8'h24; rom['h703]=8'hA0;
    rom['h704]=8'h55; rom['h705]=8'h88; rom['h706]=8'h24; rom['h707]=8'hA4;
    rom['h708]=8'h55; rom['h709]=8'h9B; rom['h70A]=8'h55; rom['h70B]=8'h42;
    rom['h70C]=8'h22; rom['h70D]=8'hA0; rom['h70E]=8'h24; rom['h70F]=8'hA4;
    rom['h710]=8'hD0; rom['h711]=8'hBA; rom['h712]=8'h56; rom['h713]=8'hA8;
    rom['h714]=8'h1A; rom['h715]=8'h18; rom['h716]=8'h56; rom['h717]=8'hC0;
    rom['h718]=8'h56; rom['h719]=8'h99; rom['h71A]=8'h7A; rom['h71B]=8'h12;
    rom['h71C]=8'h59; rom['h71D]=8'hBF; rom['h71E]=8'h59; rom['h71F]=8'hA5;
    rom['h720]=8'hC0; rom['h721]=8'h59; rom['h722]=8'hD9; rom['h723]=8'h59;
    rom['h724]=8'h5B; rom['h725]=8'h59; rom['h726]=8'h43; rom['h727]=8'h56;
    rom['h728]=8'h4C; rom['h729]=8'h24; rom['h72A]=8'h00; rom['h72B]=8'h55;
    rom['h72C]=8'hAE; rom['h72D]=8'h1A; rom['h72E]=8'h37; rom['h72F]=8'h55;
    rom['h730]=8'hEB; rom['h731]=8'h55; rom['h732]=8'hCA; rom['h733]=8'h56;
    rom['h734]=8'h52; rom['h735]=8'h24; rom['h736]=8'h01; rom['h737]=8'h59;
    rom['h738]=8'h73; rom['h739]=8'h56; rom['h73A]=8'h75; rom['h73B]=8'h20;
    rom['h73C]=8'h90; rom['h73D]=8'h55; rom['h73E]=8'hF9; rom['h73F]=8'hA2;
    rom['h740]=8'hB0; rom['h741]=8'hA3; rom['h742]=8'hB1; rom['h743]=8'h55;
    rom['h744]=8'hAE; rom['h745]=8'h1A; rom['h746]=8'h4D; rom['h747]=8'h55;
    rom['h748]=8'hEB; rom['h749]=8'h55; rom['h74A]=8'hCA; rom['h74B]=8'h56;
    rom['h74C]=8'h52; rom['h74D]=8'h56; rom['h74E]=8'h23; rom['h74F]=8'h20;
    rom['h750]=8'h90; rom['h751]=8'h28; rom['h752]=8'h00; rom['h753]=8'h2A;
    rom['h754]=8'h00; rom['h755]=8'hA4; rom['h756]=8'h1C; rom['h757]=8'h9B;
    rom['h758]=8'h56; rom['h759]=8'hF5; rom['h75A]=8'hA4; rom['h75B]=8'h1C;
    rom['h75C]=8'h8E; rom['h75D]=8'h56; rom['h75E]=8'hF5; rom['h75F]=8'hA4;
    rom['h760]=8'h1C; rom['h761]=8'h81; rom['h762]=8'h56; rom['h763]=8'hF5;
    rom['h764]=8'hA4; rom['h765]=8'h1C; rom['h766]=8'h74; rom['h767]=8'h20;
    rom['h768]=8'h90; rom['h769]=8'h55; rom['h76A]=8'h42; rom['h76B]=8'h59;
    rom['h76C]=8'h8B; rom['h76D]=8'h24; rom['h76E]=8'h7F; rom['h76F]=8'h26;
    rom['h770]=8'hFF; rom['h771]=8'h55; rom['h772]=8'hF9; rom['h773]=8'hC1;
    rom['h774]=8'h56; rom['h775]=8'h0E; rom['h776]=8'h56; rom['h777]=8'hD5;
    rom['h778]=8'h1A; rom['h779]=8'h7D; rom['h77A]=8'h68; rom['h77B]=8'h47;
    rom['h77C]=8'h76; rom['h77D]=8'h56; rom['h77E]=8'hC0; rom['h77F]=8'h56;
    rom['h780]=8'hEC; rom['h781]=8'h56; rom['h782]=8'h0E; rom['h783]=8'h56;
    rom['h784]=8'hD5; rom['h785]=8'h1A; rom['h786]=8'h8A; rom['h787]=8'h69;
    rom['h788]=8'h47; rom['h789]=8'h83; rom['h78A]=8'h56; rom['h78B]=8'hC0;
    rom['h78C]=8'h56; rom['h78D]=8'hEC; rom['h78E]=8'h56; rom['h78F]=8'h0E;
    rom['h790]=8'h56; rom['h791]=8'hD5; rom['h792]=8'h1A; rom['h793]=8'h97;
    rom['h794]=8'h6A; rom['h795]=8'h47; rom['h796]=8'h90; rom['h797]=8'h56;
    rom['h798]=8'hC0; rom['h799]=8'h56; rom['h79A]=8'hEC; rom['h79B]=8'h56;
    rom['h79C]=8'h0E; rom['h79D]=8'h56; rom['h79E]=8'hD5; rom['h79F]=8'h1A;
    rom['h7A0]=8'hA4; rom['h7A1]=8'h6B; rom['h7A2]=8'h47; rom['h7A3]=8'h9D;
    rom['h7A4]=8'h56; rom['h7A5]=8'hC0; rom['h7A6]=8'h59; rom['h7A7]=8'hBF;
    rom['h7A8]=8'hA5; rom['h7A9]=8'h14; rom['h7AA]=8'hAF; rom['h7AB]=8'h55;
    rom['h7AC]=8'hEB; rom['h7AD]=8'h55; rom['h7AE]=8'hCA; rom['h7AF]=8'hA8;
    rom['h7B0]=8'hB4; rom['h7B1]=8'hA9; rom['h7B2]=8'hB5; rom['h7B3]=8'hAA;
    rom['h7B4]=8'hB6; rom['h7B5]=8'hAB; rom['h7B6]=8'hB7; rom['h7B7]=8'h59;
    rom['h7B8]=8'h8B; rom['h7B9]=8'h55; rom['h7BA]=8'hF9; rom['h7BB]=8'h56;
    rom['h7BC]=8'h59; rom['h7BD]=8'h1A; rom['h7BE]=8'hC3; rom['h7BF]=8'h55;
    rom['h7C0]=8'hEB; rom['h7C1]=8'h55; rom['h7C2]=8'hCA; rom['h7C3]=8'h59;
    rom['h7C4]=8'hA5; rom['h7C5]=8'h59; rom['h7C6]=8'hFC; rom['h7C7]=8'hC0;
    rom['h7C8]=8'hA1; rom['h7C9]=8'hBF; rom['h7CA]=8'hA3; rom['h7CB]=8'hBD;
    rom['h7CC]=8'hF0; rom['h7CD]=8'hBC; rom['h7CE]=8'hDC; rom['h7CF]=8'hBE;
    rom['h7D0]=8'hFA; rom['h7D1]=8'hF3; rom['h7D2]=8'h21; rom['h7D3]=8'hE9;
    rom['h7D4]=8'h23; rom['h7D5]=8'hE8; rom['h7D6]=8'h61; rom['h7D7]=8'h63;
    rom['h7D8]=8'hBB; rom['h7D9]=8'hAB; rom['h7DA]=8'h14; rom['h7DB]=8'hDE;
    rom['h7DC]=8'hD1; rom['h7DD]=8'hBC; rom['h7DE]=8'h7E; rom['h7DF]=8'hD1;
    rom['h7E0]=8'hAB; rom['h7E1]=8'hF5; rom['h7E2]=8'hF3; rom['h7E3]=8'hAF;
    rom['h7E4]=8'hB1; rom['h7E5]=8'hAD; rom['h7E6]=8'hB3; rom['h7E7]=8'hAC;
    rom['h7E8]=8'h14; rom['h7E9]=8'hEB; rom['h7EA]=8'hC1; rom['h7EB]=8'hC0;
    rom['h7EC]=8'h59; rom['h7ED]=8'h73; rom['h7EE]=8'h59; rom['h7EF]=8'h5B;
    rom['h7F0]=8'h22; rom['h7F1]=8'h00; rom['h7F2]=8'h47; rom['h7F3]=8'hF8;
    rom['h7F4]=8'h59; rom['h7F5]=8'h73; rom['h7F6]=8'h59; rom['h7F7]=8'h5B;
    rom['h7F8]=8'h59; rom['h7F9]=8'h43; rom['h7FA]=8'hA2; rom['h7FB]=8'hB4;
    rom['h7FC]=8'hA3; rom['h7FD]=8'hB5; rom['h7FE]=8'h59; rom['h7FF]=8'h06;
    rom['h800]=8'h5D; rom['h801]=8'hF5; rom['h802]=8'h14; rom['h803]=8'h0E;
    rom['h804]=8'h5D; rom['h805]=8'hDD; rom['h806]=8'h14; rom['h807]=8'h0E;
    rom['h808]=8'h5D; rom['h809]=8'h28; rom['h80A]=8'h55; rom['h80B]=8'hCA;
    rom['h80C]=8'h47; rom['h80D]=8'hFE; rom['h80E]=8'h24; rom['h80F]=8'h00;
    rom['h810]=8'h5D; rom['h811]=8'hDD; rom['h812]=8'h14; rom['h813]=8'h16;
    rom['h814]=8'h55; rom['h815]=8'hCA; rom['h816]=8'h59; rom['h817]=8'h8B;
    rom['h818]=8'h59; rom['h819]=8'hA5; rom['h81A]=8'h59; rom['h81B]=8'hBF;
    rom['h81C]=8'hC0; rom['h81D]=8'h59; rom['h81E]=8'h43; rom['h81F]=8'h59;
    rom['h820]=8'hD9; rom['h821]=8'h59; rom['h822]=8'h5B; rom['h823]=8'h59;
    rom['h824]=8'h73; rom['h825]=8'hA2; rom['h826]=8'hB0; rom['h827]=8'hA3;
    rom['h828]=8'hB1; rom['h829]=8'h22; rom['h82A]=8'h90; rom['h82B]=8'h59;
    rom['h82C]=8'hD9; rom['h82D]=8'h2E; rom['h82E]=8'h7C; rom['h82F]=8'hD1;
    rom['h830]=8'h2F; rom['h831]=8'hE0; rom['h832]=8'h55; rom['h833]=8'hAE;
    rom['h834]=8'h1A; rom['h835]=8'h3E; rom['h836]=8'h55; rom['h837]=8'hEB;
    rom['h838]=8'h55; rom['h839]=8'hCA; rom['h83A]=8'h22; rom['h83B]=8'h2D;
    rom['h83C]=8'h5D; rom['h83D]=8'h28; rom['h83E]=8'h22; rom['h83F]=8'hAC;
    rom['h840]=8'h24; rom['h841]=8'h27; rom['h842]=8'h26; rom['h843]=8'h10;
    rom['h844]=8'h56; rom['h845]=8'h0E; rom['h846]=8'h57; rom['h847]=8'h21;
    rom['h848]=8'h58; rom['h849]=8'hC3; rom['h84A]=8'h22; rom['h84B]=8'h90;
    rom['h84C]=8'h55; rom['h84D]=8'h4F; rom['h84E]=8'h22; rom['h84F]=8'hAC;
    rom['h850]=8'h24; rom['h851]=8'h03; rom['h852]=8'h26; rom['h853]=8'hE8;
    rom['h854]=8'h56; rom['h855]=8'h0E; rom['h856]=8'h57; rom['h857]=8'h21;
    rom['h858]=8'h58; rom['h859]=8'hC3; rom['h85A]=8'h22; rom['h85B]=8'h90;
    rom['h85C]=8'h55; rom['h85D]=8'h4F; rom['h85E]=8'h22; rom['h85F]=8'hAC;
    rom['h860]=8'h24; rom['h861]=8'h00; rom['h862]=8'h26; rom['h863]=8'h64;
    rom['h864]=8'h56; rom['h865]=8'h0E; rom['h866]=8'h57; rom['h867]=8'h21;
    rom['h868]=8'h58; rom['h869]=8'hC3; rom['h86A]=8'h22; rom['h86B]=8'h90;
    rom['h86C]=8'h55; rom['h86D]=8'h4F; rom['h86E]=8'h22; rom['h86F]=8'hAC;
    rom['h870]=8'h24; rom['h871]=8'h00; rom['h872]=8'h26; rom['h873]=8'h0A;
    rom['h874]=8'h56; rom['h875]=8'h0E; rom['h876]=8'h57; rom['h877]=8'h21;
    rom['h878]=8'h58; rom['h879]=8'hC3; rom['h87A]=8'h20; rom['h87B]=8'h90;
    rom['h87C]=8'h21; rom['h87D]=8'hE9; rom['h87E]=8'h5D; rom['h87F]=8'h48;
    rom['h880]=8'h22; rom['h881]=8'h90; rom['h882]=8'h59; rom['h883]=8'hFC;
    rom['h884]=8'h59; rom['h885]=8'hBF; rom['h886]=8'h59; rom['h887]=8'hA5;
    rom['h888]=8'h59; rom['h889]=8'hFC; rom['h88A]=8'h59; rom['h88B]=8'h8B;
    rom['h88C]=8'hC0; rom['h88D]=8'h59; rom['h88E]=8'h5B; rom['h88F]=8'h59;
    rom['h890]=8'h73; rom['h891]=8'hA6; rom['h892]=8'hB4; rom['h893]=8'hA7;
    rom['h894]=8'hB5; rom['h895]=8'h59; rom['h896]=8'h73; rom['h897]=8'h56;
    rom['h898]=8'h23; rom['h899]=8'hA4; rom['h89A]=8'h5D; rom['h89B]=8'h48;
    rom['h89C]=8'hA5; rom['h89D]=8'h5D; rom['h89E]=8'h48; rom['h89F]=8'hA6;
    rom['h8A0]=8'h5D; rom['h8A1]=8'h48; rom['h8A2]=8'hA7; rom['h8A3]=8'h5D;
    rom['h8A4]=8'h48; rom['h8A5]=8'h59; rom['h8A6]=8'hBF; rom['h8A7]=8'hA4;
    rom['h8A8]=8'hB6; rom['h8A9]=8'hA5; rom['h8AA]=8'hB7; rom['h8AB]=8'h59;
    rom['h8AC]=8'hBF; rom['h8AD]=8'h59; rom['h8AE]=8'hA5; rom['h8AF]=8'hC0;
    rom['h8B0]=8'h59; rom['h8B1]=8'h43; rom['h8B2]=8'h59; rom['h8B3]=8'h5B;
    rom['h8B4]=8'hA2; rom['h8B5]=8'hB0; rom['h8B6]=8'hA3; rom['h8B7]=8'hB1;
    rom['h8B8]=8'hA0; rom['h8B9]=8'h5D; rom['h8BA]=8'h48; rom['h8BB]=8'hA1;
    rom['h8BC]=8'h5D; rom['h8BD]=8'h48; rom['h8BE]=8'h59; rom['h8BF]=8'hA5;
    rom['h8C0]=8'h59; rom['h8C1]=8'h8B; rom['h8C2]=8'hC0; rom['h8C3]=8'h21;
    rom['h8C4]=8'hE9; rom['h8C5]=8'h1C; rom['h8C6]=8'hCE; rom['h8C7]=8'h2E;
    rom['h8C8]=8'h7C; rom['h8C9]=8'h2F; rom['h8CA]=8'hE9; rom['h8CB]=8'h14;
    rom['h8CC]=8'hCE; rom['h8CD]=8'hC1; rom['h8CE]=8'h5D; rom['h8CF]=8'h48;
    rom['h8D0]=8'h2E; rom['h8D1]=8'h7C; rom['h8D2]=8'hF0; rom['h8D3]=8'h2F;
    rom['h8D4]=8'hE0; rom['h8D5]=8'hC0; rom['h8D6]=8'h21; rom['h8D7]=8'hA3;
    rom['h8D8]=8'hE3; rom['h8D9]=8'hA2; rom['h8DA]=8'hE3; rom['h8DB]=8'hC0;
    rom['h8DC]=8'h2D; rom['h8DD]=8'hAF; rom['h8DE]=8'hE3; rom['h8DF]=8'hAE;
    rom['h8E0]=8'hE3; rom['h8E1]=8'hC0; rom['h8E2]=8'h2C; rom['h8E3]=8'hFE;
    rom['h8E4]=8'h2E; rom['h8E5]=8'h32; rom['h8E6]=8'h58; rom['h8E7]=8'hDC;
    rom['h8E8]=8'h6D; rom['h8E9]=8'h2E; rom['h8EA]=8'hC0; rom['h8EB]=8'h58;
    rom['h8EC]=8'hDC; rom['h8ED]=8'hC0; rom['h8EE]=8'h2E; rom['h8EF]=8'h00;
    rom['h8F0]=8'h2F; rom['h8F1]=8'hE1; rom['h8F2]=8'hC0; rom['h8F3]=8'h20;
    rom['h8F4]=8'h40; rom['h8F5]=8'h5E; rom['h8F6]=8'h00; rom['h8F7]=8'h5D;
    rom['h8F8]=8'h00; rom['h8F9]=8'h5D; rom['h8FA]=8'h28; rom['h8FB]=8'h5D;
    rom['h8FC]=8'hB7; rom['h8FD]=8'hA3; rom['h8FE]=8'h58; rom['h8FF]=8'hEE;
    rom['h900]=8'h58; rom['h901]=8'hE2; rom['h902]=8'h5D; rom['h903]=8'h5C;
    rom['h904]=8'h40; rom['h905]=8'h1B; rom['h906]=8'hA0; rom['h907]=8'hBC;
    rom['h908]=8'hA1; rom['h909]=8'hBD; rom['h90A]=8'h2D; rom['h90B]=8'hE9;
    rom['h90C]=8'h2E; rom['h90D]=8'h00; rom['h90E]=8'h2F; rom['h90F]=8'hE1;
    rom['h910]=8'h6D; rom['h911]=8'h2D; rom['h912]=8'hE9; rom['h913]=8'hB1;
    rom['h914]=8'h6D; rom['h915]=8'h2D; rom['h916]=8'hE9; rom['h917]=8'hB0;
    rom['h918]=8'h5F; rom['h919]=8'hFE; rom['h91A]=8'hAC; rom['h91B]=8'hB0;
    rom['h91C]=8'hAD; rom['h91D]=8'hF8; rom['h91E]=8'hF8; rom['h91F]=8'hB1;
    rom['h920]=8'hC0; rom['h921]=8'h21; rom['h922]=8'hE9; rom['h923]=8'h2E;
    rom['h924]=8'h00; rom['h925]=8'h2F; rom['h926]=8'hE1; rom['h927]=8'h61;
    rom['h928]=8'h21; rom['h929]=8'hE9; rom['h92A]=8'hBD; rom['h92B]=8'h61;
    rom['h92C]=8'h21; rom['h92D]=8'hE9; rom['h92E]=8'hBC; rom['h92F]=8'h2D;
    rom['h930]=8'hA3; rom['h931]=8'hE3; rom['h932]=8'hA2; rom['h933]=8'hE3;
    rom['h934]=8'hA1; rom['h935]=8'hF8; rom['h936]=8'hF8; rom['h937]=8'hB1;
    rom['h938]=8'hC0; rom['h939]=8'h20; rom['h93A]=8'hFC; rom['h93B]=8'h22;
    rom['h93C]=8'h00; rom['h93D]=8'h21; rom['h93E]=8'hA2; rom['h93F]=8'hE4;
    rom['h940]=8'hA3; rom['h941]=8'hE5; rom['h942]=8'hC0; rom['h943]=8'hD2;
    rom['h944]=8'hBC; rom['h945]=8'h2E; rom['h946]=8'hFC; rom['h947]=8'h2F;
    rom['h948]=8'hED; rom['h949]=8'hF1; rom['h94A]=8'h9C; rom['h94B]=8'hE5;
    rom['h94C]=8'hBF; rom['h94D]=8'hEC; rom['h94E]=8'h12; rom['h94F]=8'h51;
    rom['h950]=8'hF8; rom['h951]=8'hE4; rom['h952]=8'hBE; rom['h953]=8'h2F;
    rom['h954]=8'hA1; rom['h955]=8'hE0; rom['h956]=8'h6F; rom['h957]=8'h2F;
    rom['h958]=8'hA0; rom['h959]=8'hE0; rom['h95A]=8'hC0; rom['h95B]=8'hD2;
    rom['h95C]=8'hBC; rom['h95D]=8'h2E; rom['h95E]=8'hFC; rom['h95F]=8'h2F;
    rom['h960]=8'hED; rom['h961]=8'hF1; rom['h962]=8'h9C; rom['h963]=8'hE5;
    rom['h964]=8'hBF; rom['h965]=8'hEC; rom['h966]=8'h12; rom['h967]=8'h69;
    rom['h968]=8'hF8; rom['h969]=8'hE4; rom['h96A]=8'hBE; rom['h96B]=8'h2F;
    rom['h96C]=8'hA3; rom['h96D]=8'hE0; rom['h96E]=8'h6F; rom['h96F]=8'h2F;
    rom['h970]=8'hA2; rom['h971]=8'hE0; rom['h972]=8'hC0; rom['h973]=8'hD2;
    rom['h974]=8'hBC; rom['h975]=8'h2E; rom['h976]=8'hFC; rom['h977]=8'h2F;
    rom['h978]=8'hED; rom['h979]=8'hF1; rom['h97A]=8'h9C; rom['h97B]=8'hE5;
    rom['h97C]=8'hBF; rom['h97D]=8'hEC; rom['h97E]=8'h12; rom['h97F]=8'h81;
    rom['h980]=8'hF8; rom['h981]=8'hE4; rom['h982]=8'hBE; rom['h983]=8'h2F;
    rom['h984]=8'hA5; rom['h985]=8'hE0; rom['h986]=8'h6F; rom['h987]=8'h2F;
    rom['h988]=8'hA4; rom['h989]=8'hE0; rom['h98A]=8'hC0; rom['h98B]=8'h2E;
    rom['h98C]=8'hFC; rom['h98D]=8'h2F; rom['h98E]=8'hEC; rom['h98F]=8'hBE;
    rom['h990]=8'hED; rom['h991]=8'hBF; rom['h992]=8'h2F; rom['h993]=8'hE9;
    rom['h994]=8'hB1; rom['h995]=8'h6F; rom['h996]=8'h2F; rom['h997]=8'hE9;
    rom['h998]=8'hB0; rom['h999]=8'h2C; rom['h99A]=8'hFC; rom['h99B]=8'h2D;
    rom['h99C]=8'h6F; rom['h99D]=8'hAF; rom['h99E]=8'hE5; rom['h99F]=8'h1C;
    rom['h9A0]=8'hA4; rom['h9A1]=8'h6E; rom['h9A2]=8'hAE; rom['h9A3]=8'hE4;
    rom['h9A4]=8'hC0; rom['h9A5]=8'h2E; rom['h9A6]=8'hFC; rom['h9A7]=8'h2F;
    rom['h9A8]=8'hEC; rom['h9A9]=8'hBE; rom['h9AA]=8'hED; rom['h9AB]=8'hBF;
    rom['h9AC]=8'h2F; rom['h9AD]=8'hE9; rom['h9AE]=8'hB3; rom['h9AF]=8'h6F;
    rom['h9B0]=8'h2F; rom['h9B1]=8'hE9; rom['h9B2]=8'hB2; rom['h9B3]=8'h2C;
    rom['h9B4]=8'hFC; rom['h9B5]=8'h2D; rom['h9B6]=8'h6F; rom['h9B7]=8'hAF;
    rom['h9B8]=8'hE5; rom['h9B9]=8'h1C; rom['h9BA]=8'hBE; rom['h9BB]=8'h6E;
    rom['h9BC]=8'hAE; rom['h9BD]=8'hE4; rom['h9BE]=8'hC0; rom['h9BF]=8'h2E;
    rom['h9C0]=8'hFC; rom['h9C1]=8'h2F; rom['h9C2]=8'hEC; rom['h9C3]=8'hBE;
    rom['h9C4]=8'hED; rom['h9C5]=8'hBF; rom['h9C6]=8'h2F; rom['h9C7]=8'hE9;
    rom['h9C8]=8'hB5; rom['h9C9]=8'h6F; rom['h9CA]=8'h2F; rom['h9CB]=8'hE9;
    rom['h9CC]=8'hB4; rom['h9CD]=8'h2C; rom['h9CE]=8'hFC; rom['h9CF]=8'h2D;
    rom['h9D0]=8'h6F; rom['h9D1]=8'hAF; rom['h9D2]=8'hE5; rom['h9D3]=8'h1C;
    rom['h9D4]=8'hD8; rom['h9D5]=8'h6E; rom['h9D6]=8'hAE; rom['h9D7]=8'hE4;
    rom['h9D8]=8'hC0; rom['h9D9]=8'hA3; rom['h9DA]=8'hBD; rom['h9DB]=8'hD4;
    rom['h9DC]=8'hBC; rom['h9DD]=8'h2E; rom['h9DE]=8'hFC; rom['h9DF]=8'h2F;
    rom['h9E0]=8'hED; rom['h9E1]=8'hF1; rom['h9E2]=8'h9C; rom['h9E3]=8'hE5;
    rom['h9E4]=8'hBF; rom['h9E5]=8'hEC; rom['h9E6]=8'h12; rom['h9E7]=8'hE9;
    rom['h9E8]=8'hF8; rom['h9E9]=8'hE4; rom['h9EA]=8'hBE; rom['h9EB]=8'hDC;
    rom['h9EC]=8'hBC; rom['h9ED]=8'h23; rom['h9EE]=8'hE9; rom['h9EF]=8'h2F;
    rom['h9F0]=8'hE0; rom['h9F1]=8'h6F; rom['h9F2]=8'hAF; rom['h9F3]=8'h1C;
    rom['h9F4]=8'hF6; rom['h9F5]=8'h6E; rom['h9F6]=8'h63; rom['h9F7]=8'h7C;
    rom['h9F8]=8'hED; rom['h9F9]=8'hAD; rom['h9FA]=8'hB3; rom['h9FB]=8'hC0;
    rom['h9FC]=8'hA3; rom['h9FD]=8'hBD; rom['h9FE]=8'h2E; rom['h9FF]=8'hFC;
    rom['hA00]=8'h2F; rom['hA01]=8'hEC; rom['hA02]=8'hBE; rom['hA03]=8'hED;
    rom['hA04]=8'hBF; rom['hA05]=8'hDC; rom['hA06]=8'hBC; rom['hA07]=8'h2F;
    rom['hA08]=8'hE9; rom['hA09]=8'h23; rom['hA0A]=8'hE0; rom['hA0B]=8'h6F;
    rom['hA0C]=8'hAF; rom['hA0D]=8'h1C; rom['hA0E]=8'h10; rom['hA0F]=8'h6E;
    rom['hA10]=8'h63; rom['hA11]=8'h7C; rom['hA12]=8'h07; rom['hA13]=8'hAD;
    rom['hA14]=8'hB3; rom['hA15]=8'h2C; rom['hA16]=8'hFC; rom['hA17]=8'h2D;
    rom['hA18]=8'hAE; rom['hA19]=8'hE4; rom['hA1A]=8'hAF; rom['hA1B]=8'hE5;
    rom['hA1C]=8'hC0; rom['hA1D]=8'h59; rom['hA1E]=8'h43; rom['hA1F]=8'h59;
    rom['hA20]=8'h5B; rom['hA21]=8'h22; rom['hA22]=8'hA0; rom['hA23]=8'h55;
    rom['hA24]=8'h62; rom['hA25]=8'h5D; rom['hA26]=8'h00; rom['hA27]=8'h5C;
    rom['hA28]=8'hEF; rom['hA29]=8'h14; rom['hA2A]=8'h31; rom['hA2B]=8'h5D;
    rom['hA2C]=8'h69; rom['hA2D]=8'h5D; rom['hA2E]=8'h6D; rom['hA2F]=8'h4A;
    rom['hA30]=8'h53; rom['hA31]=8'h2E; rom['hA32]=8'h08; rom['hA33]=8'h5D;
    rom['hA34]=8'hD0; rom['hA35]=8'h1C; rom['hA36]=8'h4B; rom['hA37]=8'h22;
    rom['hA38]=8'hA0; rom['hA39]=8'h57; rom['hA3A]=8'hC8; rom['hA3B]=8'h1C;
    rom['hA3C]=8'h3F; rom['hA3D]=8'h4A; rom['hA3E]=8'h25; rom['hA3F]=8'h55;
    rom['hA40]=8'hDA; rom['hA41]=8'h22; rom['hA42]=8'h08; rom['hA43]=8'h5D;
    rom['hA44]=8'h28; rom['hA45]=8'h5D; rom['hA46]=8'h53; rom['hA47]=8'h5D;
    rom['hA48]=8'h28; rom['hA49]=8'h4A; rom['hA4A]=8'h25; rom['hA4B]=8'h5D;
    rom['hA4C]=8'h28; rom['hA4D]=8'h59; rom['hA4E]=8'h21; rom['hA4F]=8'h55;
    rom['hA50]=8'hCA; rom['hA51]=8'h4A; rom['hA52]=8'h25; rom['hA53]=8'h22;
    rom['hA54]=8'h00; rom['hA55]=8'h59; rom['hA56]=8'h21; rom['hA57]=8'h55;
    rom['hA58]=8'hCA; rom['hA59]=8'h59; rom['hA5A]=8'h21; rom['hA5B]=8'h22;
    rom['hA5C]=8'hA0; rom['hA5D]=8'h55; rom['hA5E]=8'h4F; rom['hA5F]=8'h59;
    rom['hA60]=8'hA5; rom['hA61]=8'h59; rom['hA62]=8'h8B; rom['hA63]=8'hC0;
    rom['hA64]=8'h59; rom['hA65]=8'h43; rom['hA66]=8'h59; rom['hA67]=8'h5B;
    rom['hA68]=8'hA0; rom['hA69]=8'hB4; rom['hA6A]=8'hA1; rom['hA6B]=8'hB5;
    rom['hA6C]=8'hA2; rom['hA6D]=8'hB0; rom['hA6E]=8'hA3; rom['hA6F]=8'hB1;
    rom['hA70]=8'h55; rom['hA71]=8'h42; rom['hA72]=8'h20; rom['hA73]=8'hA0;
    rom['hA74]=8'h55; rom['hA75]=8'h42; rom['hA76]=8'hA4; rom['hA77]=8'hB0;
    rom['hA78]=8'hA5; rom['hA79]=8'hB1; rom['hA7A]=8'h59; rom['hA7B]=8'h06;
    rom['hA7C]=8'h2E; rom['hA7D]=8'h30; rom['hA7E]=8'h5D; rom['hA7F]=8'hD0;
    rom['hA80]=8'h1C; rom['hA81]=8'h84; rom['hA82]=8'h4A; rom['hA83]=8'hBF;
    rom['hA84]=8'h5D; rom['hA85]=8'hB7; rom['hA86]=8'h20; rom['hA87]=8'hA4;
    rom['hA88]=8'h56; rom['hA89]=8'h38; rom['hA8A]=8'h20; rom['hA8B]=8'hA0;
    rom['hA8C]=8'h22; rom['hA8D]=8'hA0; rom['hA8E]=8'h55; rom['hA8F]=8'hB9;
    rom['hA90]=8'h14; rom['hA91]=8'h9E; rom['hA92]=8'h22; rom['hA93]=8'hA8;
    rom['hA94]=8'h55; rom['hA95]=8'h62; rom['hA96]=8'h56; rom['hA97]=8'h8A;
    rom['hA98]=8'h56; rom['hA99]=8'h8A; rom['hA9A]=8'h56; rom['hA9B]=8'hC0;
    rom['hA9C]=8'h56; rom['hA9D]=8'h8A; rom['hA9E]=8'h22; rom['hA9F]=8'hA4;
    rom['hAA0]=8'h56; rom['hAA1]=8'hC0; rom['hAA2]=8'hA4; rom['hAA3]=8'hB0;
    rom['hAA4]=8'hA5; rom['hAA5]=8'hB1; rom['hAA6]=8'h55; rom['hAA7]=8'hCA;
    rom['hAA8]=8'h59; rom['hAA9]=8'h06; rom['hAAA]=8'h5D; rom['hAAB]=8'h8C;
    rom['hAAC]=8'h14; rom['hAAD]=8'hB0; rom['hAAE]=8'h4A; rom['hAAF]=8'h84;
    rom['hAB0]=8'h59; rom['hAB1]=8'hA5; rom['hAB2]=8'h20; rom['hAB3]=8'hA0;
    rom['hAB4]=8'h55; rom['hAB5]=8'h62; rom['hAB6]=8'h59; rom['hAB7]=8'h8B;
    rom['hAB8]=8'hC0; rom['hAB9]=8'h20; rom['hABA]=8'hA0; rom['hABB]=8'h55;
    rom['hABC]=8'hF9; rom['hABD]=8'h4A; rom['hABE]=8'hB0; rom['hABF]=8'h24;
    rom['hAC0]=8'h00; rom['hAC1]=8'h26; rom['hAC2]=8'h00; rom['hAC3]=8'h55;
    rom['hAC4]=8'hCA; rom['hAC5]=8'h59; rom['hAC6]=8'h06; rom['hAC7]=8'h50;
    rom['hAC8]=8'hA6; rom['hAC9]=8'h14; rom['hACA]=8'hB9; rom['hACB]=8'h5D;
    rom['hACC]=8'hB7; rom['hACD]=8'h56; rom['hACE]=8'hF5; rom['hACF]=8'hA3;
    rom['hAD0]=8'hB7; rom['hAD1]=8'h4A; rom['hAD2]=8'hC3; rom['hAD3]=8'h20;
    rom['hAD4]=8'h4E; rom['hAD5]=8'h5E; rom['hAD6]=8'h00; rom['hAD7]=8'hF0;
    rom['hAD8]=8'hB4; rom['hAD9]=8'h5D; rom['hADA]=8'h00; rom['hADB]=8'h5D;
    rom['hADC]=8'h28; rom['hADD]=8'h5D; rom['hADE]=8'hB7; rom['hADF]=8'hA3;
    rom['hAE0]=8'hB5; rom['hAE1]=8'h5D; rom['hAE2]=8'h00; rom['hAE3]=8'h5D;
    rom['hAE4]=8'h28; rom['hAE5]=8'h5D; rom['hAE6]=8'hB7; rom['hAE7]=8'hA3;
    rom['hAE8]=8'hB6; rom['hAE9]=8'hF0; rom['hAEA]=8'hB7; rom['hAEB]=8'h22;
    rom['hAEC]=8'hA0; rom['hAED]=8'h56; rom['hAEE]=8'h0E; rom['hAEF]=8'h5D;
    rom['hAF0]=8'h00; rom['hAF1]=8'h5D; rom['hAF2]=8'h28; rom['hAF3]=8'h5D;
    rom['hAF4]=8'hB7; rom['hAF5]=8'hA3; rom['hAF6]=8'hF4; rom['hAF7]=8'hBB;
    rom['hAF8]=8'h00; rom['hAF9]=8'h00; rom['hAFA]=8'h00; rom['hAFB]=8'h00;
    rom['hAFC]=8'h00; rom['hAFD]=8'h00; rom['hAFE]=8'h00; rom['hAFF]=8'h00;
    rom['hB00]=8'h5D; rom['hB01]=8'h5C; rom['hB02]=8'h22; rom['hB03]=8'hA0;
    rom['hB04]=8'h58; rom['hB05]=8'h8D; rom['hB06]=8'h22; rom['hB07]=8'h3A;
    rom['hB08]=8'h5D; rom['hB09]=8'h28; rom['hB0A]=8'hD0; rom['hB0B]=8'hBA;
    rom['hB0C]=8'h20; rom['hB0D]=8'hA0; rom['hB0E]=8'h59; rom['hB0F]=8'h06;
    rom['hB10]=8'h58; rom['hB11]=8'hB0; rom['hB12]=8'h55; rom['hB13]=8'hCA;
    rom['hB14]=8'h7A; rom['hB15]=8'h0C; rom['hB16]=8'h7B; rom['hB17]=8'h00;
    rom['hB18]=8'h5D; rom['hB19]=8'h5C; rom['hB1A]=8'h40; rom['hB1B]=8'h1B;
    rom['hB1C]=8'h20; rom['hB1D]=8'h4E; rom['hB1E]=8'h5E; rom['hB1F]=8'h00;
    rom['hB20]=8'hF0; rom['hB21]=8'hB4; rom['hB22]=8'h5D; rom['hB23]=8'h00;
    rom['hB24]=8'h5D; rom['hB25]=8'h28; rom['hB26]=8'h5D; rom['hB27]=8'hB7;
    rom['hB28]=8'hA3; rom['hB29]=8'hB5; rom['hB2A]=8'h5D; rom['hB2B]=8'h00;
    rom['hB2C]=8'h5D; rom['hB2D]=8'h28; rom['hB2E]=8'h5D; rom['hB2F]=8'hB7;
    rom['hB30]=8'hA3; rom['hB31]=8'hB6; rom['hB32]=8'h5D; rom['hB33]=8'h00;
    rom['hB34]=8'h5D; rom['hB35]=8'h28; rom['hB36]=8'h5D; rom['hB37]=8'hB7;
    rom['hB38]=8'hA3; rom['hB39]=8'hB7; rom['hB3A]=8'h22; rom['hB3B]=8'hA0;
    rom['hB3C]=8'h56; rom['hB3D]=8'h0E; rom['hB3E]=8'h5D; rom['hB3F]=8'h5C;
    rom['hB40]=8'h22; rom['hB41]=8'hA0; rom['hB42]=8'h58; rom['hB43]=8'h8D;
    rom['hB44]=8'h22; rom['hB45]=8'h3A; rom['hB46]=8'h5D; rom['hB47]=8'h28;
    rom['hB48]=8'h5D; rom['hB49]=8'h00; rom['hB4A]=8'h5C; rom['hB4B]=8'hEF;
    rom['hB4C]=8'h1C; rom['hB4D]=8'h64; rom['hB4E]=8'h5D; rom['hB4F]=8'h28;
    rom['hB50]=8'h5D; rom['hB51]=8'hB7; rom['hB52]=8'hA3; rom['hB53]=8'hB4;
    rom['hB54]=8'h5D; rom['hB55]=8'h00; rom['hB56]=8'h5D; rom['hB57]=8'h28;
    rom['hB58]=8'h5D; rom['hB59]=8'hB7; rom['hB5A]=8'hA4; rom['hB5B]=8'hB2;
    rom['hB5C]=8'h20; rom['hB5D]=8'hA0; rom['hB5E]=8'h59; rom['hB5F]=8'h21;
    rom['hB60]=8'h55; rom['hB61]=8'hCA; rom['hB62]=8'h4B; rom['hB63]=8'h3E;
    rom['hB64]=8'h5D; rom['hB65]=8'h5C; rom['hB66]=8'h40; rom['hB67]=8'h1B;
    rom['hB68]=8'hFF; rom['hB69]=8'hFF; rom['hB6A]=8'hFF; rom['hB6B]=8'hFF;
    rom['hB6C]=8'hFF; rom['hB6D]=8'hFF; rom['hB6E]=8'hFF; rom['hB6F]=8'hFF;
    rom['hB70]=8'hFF; rom['hB71]=8'hFF; rom['hB72]=8'hFF; rom['hB73]=8'hFF;
    rom['hB74]=8'hFF; rom['hB75]=8'hFF; rom['hB76]=8'hFF; rom['hB77]=8'hFF;
    rom['hB78]=8'hFF; rom['hB79]=8'hFF; rom['hB7A]=8'hFF; rom['hB7B]=8'hFF;
    rom['hB7C]=8'hFF; rom['hB7D]=8'hFF; rom['hB7E]=8'hFF; rom['hB7F]=8'hFF;
    rom['hB80]=8'hFF; rom['hB81]=8'hFF; rom['hB82]=8'hFF; rom['hB83]=8'hFF;
    rom['hB84]=8'hFF; rom['hB85]=8'hFF; rom['hB86]=8'hFF; rom['hB87]=8'hFF;
    rom['hB88]=8'hFF; rom['hB89]=8'hFF; rom['hB8A]=8'hFF; rom['hB8B]=8'hFF;
    rom['hB8C]=8'hFF; rom['hB8D]=8'hFF; rom['hB8E]=8'hFF; rom['hB8F]=8'hFF;
    rom['hB90]=8'hFF; rom['hB91]=8'hFF; rom['hB92]=8'hFF; rom['hB93]=8'hFF;
    rom['hB94]=8'hFF; rom['hB95]=8'hFF; rom['hB96]=8'hFF; rom['hB97]=8'hFF;
    rom['hB98]=8'hFF; rom['hB99]=8'hFF; rom['hB9A]=8'hFF; rom['hB9B]=8'hFF;
    rom['hB9C]=8'hFF; rom['hB9D]=8'hFF; rom['hB9E]=8'hFF; rom['hB9F]=8'hFF;
    rom['hBA0]=8'hFF; rom['hBA1]=8'hFF; rom['hBA2]=8'hFF; rom['hBA3]=8'hFF;
    rom['hBA4]=8'hFF; rom['hBA5]=8'hFF; rom['hBA6]=8'hFF; rom['hBA7]=8'hFF;
    rom['hBA8]=8'hFF; rom['hBA9]=8'hFF; rom['hBAA]=8'hFF; rom['hBAB]=8'hFF;
    rom['hBAC]=8'hFF; rom['hBAD]=8'hFF; rom['hBAE]=8'hFF; rom['hBAF]=8'hFF;
    rom['hBB0]=8'hFF; rom['hBB1]=8'hFF; rom['hBB2]=8'hFF; rom['hBB3]=8'hFF;
    rom['hBB4]=8'hFF; rom['hBB5]=8'hFF; rom['hBB6]=8'hFF; rom['hBB7]=8'hFF;
    rom['hBB8]=8'hFF; rom['hBB9]=8'hFF; rom['hBBA]=8'hFF; rom['hBBB]=8'hFF;
    rom['hBBC]=8'hFF; rom['hBBD]=8'hFF; rom['hBBE]=8'hFF; rom['hBBF]=8'hFF;
    rom['hBC0]=8'hFF; rom['hBC1]=8'hFF; rom['hBC2]=8'hFF; rom['hBC3]=8'hFF;
    rom['hBC4]=8'hFF; rom['hBC5]=8'hFF; rom['hBC6]=8'hFF; rom['hBC7]=8'hFF;
    rom['hBC8]=8'hFF; rom['hBC9]=8'hFF; rom['hBCA]=8'hFF; rom['hBCB]=8'hFF;
    rom['hBCC]=8'hFF; rom['hBCD]=8'hFF; rom['hBCE]=8'hFF; rom['hBCF]=8'hFF;
    rom['hBD0]=8'hA5; rom['hBD1]=8'h1C; rom['hBD2]=8'hDC; rom['hBD3]=8'hA4;
    rom['hBD4]=8'h1C; rom['hBD5]=8'hDC; rom['hBD6]=8'h20; rom['hBD7]=8'h78;
    rom['hBD8]=8'h22; rom['hBD9]=8'hB0; rom['hBDA]=8'h41; rom['hBDB]=8'h16;
    rom['hBDC]=8'h35; rom['hBDD]=8'h42; rom['hBDE]=8'hC7; rom['hBDF]=8'h43;
    rom['hBE0]=8'hAE; rom['hBE1]=8'h43; rom['hBE2]=8'hD6; rom['hBE3]=8'h44;
    rom['hBE4]=8'h66; rom['hBE5]=8'h44; rom['hBE6]=8'h78; rom['hBE7]=8'h43;
    rom['hBE8]=8'h5C; rom['hBE9]=8'h44; rom['hBEA]=8'hFC; rom['hBEB]=8'hFF;
    rom['hBEC]=8'hFF; rom['hBED]=8'hFF; rom['hBEE]=8'hFF; rom['hBEF]=8'hFF;
    rom['hBF0]=8'hFF; rom['hBF1]=8'hFF; rom['hBF2]=8'hFF; rom['hBF3]=8'hFF;
    rom['hBF4]=8'hFF; rom['hBF5]=8'hFF; rom['hBF6]=8'hFF; rom['hBF7]=8'hFF;
    rom['hBF8]=8'hFF; rom['hBF9]=8'hFF; rom['hBFA]=8'hFF; rom['hBFB]=8'hFF;
    rom['hBFC]=8'hFF; rom['hBFD]=8'hFF; rom['hBFE]=8'hFF; rom['hBFF]=8'hFF;
    rom['hC00]=8'h5D; rom['hC01]=8'h5C; rom['hC02]=8'h5F; rom['hC03]=8'h00;
    rom['hC04]=8'h40; rom['hC05]=8'h1B; rom['hC06]=8'hDC; rom['hC07]=8'hB4;
    rom['hC08]=8'hD0; rom['hC09]=8'hB7; rom['hC0A]=8'hF0; rom['hC0B]=8'hD4;
    rom['hC0C]=8'h84; rom['hC0D]=8'hF1; rom['hC0E]=8'h8B; rom['hC0F]=8'hB6;
    rom['hC10]=8'h27; rom['hC11]=8'hE9; rom['hC12]=8'h5D; rom['hC13]=8'h48;
    rom['hC14]=8'h77; rom['hC15]=8'h0A; rom['hC16]=8'h22; rom['hC17]=8'h3A;
    rom['hC18]=8'h5D; rom['hC19]=8'h28; rom['hC1A]=8'h27; rom['hC1B]=8'hEC;
    rom['hC1C]=8'h5D; rom['hC1D]=8'h48; rom['hC1E]=8'h27; rom['hC1F]=8'hED;
    rom['hC20]=8'h5D; rom['hC21]=8'h48; rom['hC22]=8'h27; rom['hC23]=8'hEE;
    rom['hC24]=8'h5D; rom['hC25]=8'h48; rom['hC26]=8'h27; rom['hC27]=8'hEF;
    rom['hC28]=8'h5D; rom['hC29]=8'h48; rom['hC2A]=8'h5D; rom['hC2B]=8'h5C;
    rom['hC2C]=8'h74; rom['hC2D]=8'h08; rom['hC2E]=8'h40; rom['hC2F]=8'h1B;
    rom['hC30]=8'hDC; rom['hC31]=8'hB4; rom['hC32]=8'hD0; rom['hC33]=8'hB7;
    rom['hC34]=8'hF0; rom['hC35]=8'hD4; rom['hC36]=8'h84; rom['hC37]=8'hF1;
    rom['hC38]=8'h8B; rom['hC39]=8'hB6; rom['hC3A]=8'h5D; rom['hC3B]=8'h00;
    rom['hC3C]=8'h5D; rom['hC3D]=8'hB7; rom['hC3E]=8'h27; rom['hC3F]=8'hA3;
    rom['hC40]=8'hE0; rom['hC41]=8'h5D; rom['hC42]=8'h48; rom['hC43]=8'h77;
    rom['hC44]=8'h34; rom['hC45]=8'h22; rom['hC46]=8'h3A; rom['hC47]=8'h5D;
    rom['hC48]=8'h28; rom['hC49]=8'h5D; rom['hC4A]=8'h00; rom['hC4B]=8'h5D;
    rom['hC4C]=8'hB7; rom['hC4D]=8'h27; rom['hC4E]=8'hA3; rom['hC4F]=8'hE4;
    rom['hC50]=8'h5D; rom['hC51]=8'h48; rom['hC52]=8'h5D; rom['hC53]=8'h00;
    rom['hC54]=8'h5D; rom['hC55]=8'hB7; rom['hC56]=8'h27; rom['hC57]=8'hA3;
    rom['hC58]=8'hE5; rom['hC59]=8'h5D; rom['hC5A]=8'h48; rom['hC5B]=8'h5D;
    rom['hC5C]=8'h00; rom['hC5D]=8'h5D; rom['hC5E]=8'hB7; rom['hC5F]=8'h27;
    rom['hC60]=8'hA3; rom['hC61]=8'hE6; rom['hC62]=8'h5D; rom['hC63]=8'h48;
    rom['hC64]=8'h5D; rom['hC65]=8'h00; rom['hC66]=8'h5D; rom['hC67]=8'hB7;
    rom['hC68]=8'h27; rom['hC69]=8'hA3; rom['hC6A]=8'hE7; rom['hC6B]=8'h5D;
    rom['hC6C]=8'h48; rom['hC6D]=8'h5D; rom['hC6E]=8'h5C; rom['hC6F]=8'h74;
    rom['hC70]=8'h32; rom['hC71]=8'h40; rom['hC72]=8'h1B; rom['hC73]=8'h20;
    rom['hC74]=8'h4E; rom['hC75]=8'h5E; rom['hC76]=8'h00; rom['hC77]=8'h5D;
    rom['hC78]=8'h00; rom['hC79]=8'h5D; rom['hC7A]=8'h28; rom['hC7B]=8'h5D;
    rom['hC7C]=8'hB7; rom['hC7D]=8'hA3; rom['hC7E]=8'hB5; rom['hC7F]=8'h5D;
    rom['hC80]=8'h5C; rom['hC81]=8'h22; rom['hC82]=8'h46; rom['hC83]=8'h5D;
    rom['hC84]=8'h28; rom['hC85]=8'hA5; rom['hC86]=8'h5D; rom['hC87]=8'h48;
    rom['hC88]=8'h22; rom['hC89]=8'h30; rom['hC8A]=8'h5D; rom['hC8B]=8'h28;
    rom['hC8C]=8'h22; rom['hC8D]=8'h3A; rom['hC8E]=8'h5D; rom['hC8F]=8'h28;
    rom['hC90]=8'hA5; rom['hC91]=8'hB0; rom['hC92]=8'hD0; rom['hC93]=8'hB1;
    rom['hC94]=8'h5D; rom['hC95]=8'h53; rom['hC96]=8'h5D; rom['hC97]=8'h00;
    rom['hC98]=8'h5D; rom['hC99]=8'h28; rom['hC9A]=8'h5D; rom['hC9B]=8'hB7;
    rom['hC9C]=8'hA3; rom['hC9D]=8'hB4; rom['hC9E]=8'h5D; rom['hC9F]=8'h00;
    rom['hCA0]=8'h5D; rom['hCA1]=8'h28; rom['hCA2]=8'h5D; rom['hCA3]=8'hB7;
    rom['hCA4]=8'hA4; rom['hCA5]=8'hB2; rom['hCA6]=8'h58; rom['hCA7]=8'hD6;
    rom['hCA8]=8'h71; rom['hCA9]=8'h94; rom['hCAA]=8'h5D; rom['hCAB]=8'h5C;
    rom['hCAC]=8'h40; rom['hCAD]=8'h1B; rom['hCAE]=8'h5D; rom['hCAF]=8'h5C;
    rom['hCB0]=8'h58; rom['hCB1]=8'hE2; rom['hCB2]=8'h20; rom['hCB3]=8'h00;
    rom['hCB4]=8'h22; rom['hCB5]=8'h46; rom['hCB6]=8'h5D; rom['hCB7]=8'h28;
    rom['hCB8]=8'hA0; rom['hCB9]=8'h5D; rom['hCBA]=8'h48; rom['hCBB]=8'h22;
    rom['hCBC]=8'h30; rom['hCBD]=8'h5D; rom['hCBE]=8'h28; rom['hCBF]=8'h22;
    rom['hCC0]=8'h3A; rom['hCC1]=8'h5D; rom['hCC2]=8'h28; rom['hCC3]=8'h5F;
    rom['hCC4]=8'hFE; rom['hCC5]=8'hA3; rom['hCC6]=8'hB5; rom['hCC7]=8'hA2;
    rom['hCC8]=8'h5D; rom['hCC9]=8'h48; rom['hCCA]=8'hA5; rom['hCCB]=8'h5D;
    rom['hCCC]=8'h48; rom['hCCD]=8'h71; rom['hCCE]=8'hC3; rom['hCCF]=8'h5D;
    rom['hCD0]=8'h5C; rom['hCD1]=8'h70; rom['hCD2]=8'hB4; rom['hCD3]=8'h40;
    rom['hCD4]=8'h1B; rom['hCD5]=8'h5D; rom['hCD6]=8'h5C; rom['hCD7]=8'h24;
    rom['hCD8]=8'h00; rom['hCD9]=8'hA5; rom['hCDA]=8'h58; rom['hCDB]=8'hEE;
    rom['hCDC]=8'h20; rom['hCDD]=8'h00; rom['hCDE]=8'h22; rom['hCDF]=8'h00;
    rom['hCE0]=8'h58; rom['hCE1]=8'hD6; rom['hCE2]=8'h71; rom['hCE3]=8'hE0;
    rom['hCE4]=8'h70; rom['hCE5]=8'hE0; rom['hCE6]=8'h58; rom['hCE7]=8'hE2;
    rom['hCE8]=8'h75; rom['hCE9]=8'hD9; rom['hCEA]=8'hF0; rom['hCEB]=8'h58;
    rom['hCEC]=8'hEE; rom['hCED]=8'h40; rom['hCEE]=8'h1B; rom['hCEF]=8'hA2;
    rom['hCF0]=8'h1C; rom['hCF1]=8'hFC; rom['hCF2]=8'hF1; rom['hCF3]=8'hDD;
    rom['hCF4]=8'h93; rom['hCF5]=8'h14; rom['hCF6]=8'hFD; rom['hCF7]=8'hF1;
    rom['hCF8]=8'hDA; rom['hCF9]=8'h93; rom['hCFA]=8'h14; rom['hCFB]=8'hFD;
    rom['hCFC]=8'hC0; rom['hCFD]=8'hC1; rom['hCFE]=8'hFF; rom['hCFF]=8'hFF;
    rom['hD00]=8'h2C; rom['hD01]=8'h0C; rom['hD02]=8'h19; rom['hD03]=8'h02;
    rom['hD04]=8'h2E; rom['hD05]=8'h0C; rom['hD06]=8'h7F; rom['hD07]=8'h06;
    rom['hD08]=8'h19; rom['hD09]=8'h0D; rom['hD0A]=8'hF1; rom['hD0B]=8'h4D;
    rom['hD0C]=8'h10; rom['hD0D]=8'hFA; rom['hD0E]=8'h00; rom['hD0F]=8'h00;
    rom['hD10]=8'hF6; rom['hD11]=8'h00; rom['hD12]=8'h7D; rom['hD13]=8'h08;
    rom['hD14]=8'hB3; rom['hD15]=8'h2C; rom['hD16]=8'h0C; rom['hD17]=8'h19;
    rom['hD18]=8'h1C; rom['hD19]=8'hF1; rom['hD1A]=8'h4D; rom['hD1B]=8'h1F;
    rom['hD1C]=8'hFA; rom['hD1D]=8'h00; rom['hD1E]=8'h00; rom['hD1F]=8'hF6;
    rom['hD20]=8'h00; rom['hD21]=8'h7D; rom['hD22]=8'h17; rom['hD23]=8'hB2;
    rom['hD24]=8'h19; rom['hD25]=8'h27; rom['hD26]=8'hC1; rom['hD27]=8'hC0;
    rom['hD28]=8'h2E; rom['hD29]=8'hC0; rom['hD2A]=8'h2F; rom['hD2B]=8'h2C;
    rom['hD2C]=8'h0B; rom['hD2D]=8'hA3; rom['hD2E]=8'hF1; rom['hD2F]=8'hF5;
    rom['hD30]=8'h00; rom['hD31]=8'h00; rom['hD32]=8'h00; rom['hD33]=8'h00;
    rom['hD34]=8'h00; rom['hD35]=8'hE1; rom['hD36]=8'hF6; rom['hD37]=8'h7D;
    rom['hD38]=8'h30; rom['hD39]=8'h2C; rom['hD3A]=8'h0B; rom['hD3B]=8'hA2;
    rom['hD3C]=8'hFA; rom['hD3D]=8'h00; rom['hD3E]=8'h00; rom['hD3F]=8'hE1;
    rom['hD40]=8'h2E; rom['hD41]=8'h0E; rom['hD42]=8'h7F; rom['hD43]=8'h42;
    rom['hD44]=8'hF6; rom['hD45]=8'h7D; rom['hD46]=8'h3F; rom['hD47]=8'hC0;
    rom['hD48]=8'h22; rom['hD49]=8'h30; rom['hD4A]=8'hF1; rom['hD4B]=8'hFB;
    rom['hD4C]=8'h1A; rom['hD4D]=8'h50; rom['hD4E]=8'h62; rom['hD4F]=8'hF2;
    rom['hD50]=8'hB3; rom['hD51]=8'h4D; rom['hD52]=8'h28; rom['hD53]=8'h59;
    rom['hD54]=8'h5B; rom['hD55]=8'h22; rom['hD56]=8'h20; rom['hD57]=8'h5D;
    rom['hD58]=8'h28; rom['hD59]=8'h59; rom['hD5A]=8'hA5; rom['hD5B]=8'hC0;
    rom['hD5C]=8'h59; rom['hD5D]=8'h5B; rom['hD5E]=8'h22; rom['hD5F]=8'h0D;
    rom['hD60]=8'h5D; rom['hD61]=8'h28; rom['hD62]=8'h22; rom['hD63]=8'h0A;
    rom['hD64]=8'h5D; rom['hD65]=8'h28; rom['hD66]=8'h59; rom['hD67]=8'hA5;
    rom['hD68]=8'hC0; rom['hD69]=8'h22; rom['hD6A]=8'h0D; rom['hD6B]=8'h4D;
    rom['hD6C]=8'h28; rom['hD6D]=8'h22; rom['hD6E]=8'h0A; rom['hD6F]=8'h4D;
    rom['hD70]=8'h28; rom['hD71]=8'hD0; rom['hD72]=8'hFD; rom['hD73]=8'h2E;
    rom['hD74]=8'h40; rom['hD75]=8'h2F; rom['hD76]=8'hA2; rom['hD77]=8'hE1;
    rom['hD78]=8'hD0; rom['hD79]=8'hFD; rom['hD7A]=8'h2E; rom['hD7B]=8'h80;
    rom['hD7C]=8'h2F; rom['hD7D]=8'hA3; rom['hD7E]=8'hE1; rom['hD7F]=8'hD0;
    rom['hD80]=8'hFD; rom['hD81]=8'hC0; rom['hD82]=8'hD0; rom['hD83]=8'hFD;
    rom['hD84]=8'h2E; rom['hD85]=8'hC0; rom['hD86]=8'h2F; rom['hD87]=8'hD1;
    rom['hD88]=8'hE1; rom['hD89]=8'hD0; rom['hD8A]=8'hFD; rom['hD8B]=8'hC0;
    rom['hD8C]=8'h2E; rom['hD8D]=8'h30; rom['hD8E]=8'h5D; rom['hD8F]=8'hD0;
    rom['hD90]=8'h1A; rom['hD91]=8'h99; rom['hD92]=8'h2E; rom['hD93]=8'h3A;
    rom['hD94]=8'h5D; rom['hD95]=8'hD0; rom['hD96]=8'h12; rom['hD97]=8'h99;
    rom['hD98]=8'hC1; rom['hD99]=8'hC0; rom['hD9A]=8'h2E; rom['hD9B]=8'h41;
    rom['hD9C]=8'h5D; rom['hD9D]=8'hD0; rom['hD9E]=8'h12; rom['hD9F]=8'hA1;
    rom['hDA0]=8'hC0; rom['hDA1]=8'h2E; rom['hDA2]=8'h5B; rom['hDA3]=8'h5D;
    rom['hDA4]=8'hD0; rom['hDA5]=8'h12; rom['hDA6]=8'hA8; rom['hDA7]=8'hC1;
    rom['hDA8]=8'h2E; rom['hDA9]=8'h61; rom['hDAA]=8'h5D; rom['hDAB]=8'hD0;
    rom['hDAC]=8'h12; rom['hDAD]=8'hAF; rom['hDAE]=8'hC0; rom['hDAF]=8'h2E;
    rom['hDB0]=8'h7B; rom['hDB1]=8'h5D; rom['hDB2]=8'hD0; rom['hDB3]=8'h12;
    rom['hDB4]=8'hB6; rom['hDB5]=8'hC1; rom['hDB6]=8'hC0; rom['hDB7]=8'hF0;
    rom['hDB8]=8'hD3; rom['hDB9]=8'h92; rom['hDBA]=8'h14; rom['hDBB]=8'hC0;
    rom['hDBC]=8'hF0; rom['hDBD]=8'hD9; rom['hDBE]=8'h83; rom['hDBF]=8'hB3;
    rom['hDC0]=8'hF0; rom['hDC1]=8'hB2; rom['hDC2]=8'hC0; rom['hDC3]=8'hF0;
    rom['hDC4]=8'hA0; rom['hDC5]=8'h92; rom['hDC6]=8'h14; rom['hDC7]=8'hC9;
    rom['hDC8]=8'hC1; rom['hDC9]=8'hF0; rom['hDCA]=8'hA1; rom['hDCB]=8'h93;
    rom['hDCC]=8'h14; rom['hDCD]=8'hCF; rom['hDCE]=8'hC1; rom['hDCF]=8'hC0;
    rom['hDD0]=8'hF0; rom['hDD1]=8'hA2; rom['hDD2]=8'h9E; rom['hDD3]=8'h14;
    rom['hDD4]=8'hD6; rom['hDD5]=8'hC1; rom['hDD6]=8'hF0; rom['hDD7]=8'hA3;
    rom['hDD8]=8'h9F; rom['hDD9]=8'h14; rom['hDDA]=8'hDC; rom['hDDB]=8'hC1;
    rom['hDDC]=8'hC0; rom['hDDD]=8'hA2; rom['hDDE]=8'hF1; rom['hDDF]=8'h94;
    rom['hDE0]=8'h1C; rom['hDE1]=8'hE8; rom['hDE2]=8'hA3; rom['hDE3]=8'hF1;
    rom['hDE4]=8'h95; rom['hDE5]=8'h1C; rom['hDE6]=8'hE8; rom['hDE7]=8'hC0;
    rom['hDE8]=8'hC1; rom['hDE9]=8'hA4; rom['hDEA]=8'hF1; rom['hDEB]=8'h9E;
    rom['hDEC]=8'h1C; rom['hDED]=8'hF4; rom['hDEE]=8'hA5; rom['hDEF]=8'hF1;
    rom['hDF0]=8'h9F; rom['hDF1]=8'h1C; rom['hDF2]=8'hF4; rom['hDF3]=8'hC0;
    rom['hDF4]=8'hC1; rom['hDF5]=8'hA3; rom['hDF6]=8'h1C; rom['hDF7]=8'hFC;
    rom['hDF8]=8'hA2; rom['hDF9]=8'h1C; rom['hDFA]=8'hFC; rom['hDFB]=8'hC0;
    rom['hDFC]=8'hC1; rom['hDFD]=8'hFF; rom['hDFE]=8'hFF; rom['hDFF]=8'hFF;
    rom['hE00]=8'h59; rom['hE01]=8'h43; rom['hE02]=8'h59; rom['hE03]=8'h5B;
    rom['hE04]=8'h32; rom['hE05]=8'hA2; rom['hE06]=8'h1C; rom['hE07]=8'h0B;
    rom['hE08]=8'hA3; rom['hE09]=8'h14; rom['hE0A]=8'h12; rom['hE0B]=8'h5D;
    rom['hE0C]=8'h28; rom['hE0D]=8'h71; rom['hE0E]=8'h04; rom['hE0F]=8'h60;
    rom['hE10]=8'h4E; rom['hE11]=8'h04; rom['hE12]=8'h59; rom['hE13]=8'hA5;
    rom['hE14]=8'h59; rom['hE15]=8'h8B; rom['hE16]=8'hC0; rom['hE17]=8'h0D;
    rom['hE18]=8'h49; rom['hE19]=8'h6E; rom['hE1A]=8'h74; rom['hE1B]=8'h65;
    rom['hE1C]=8'h6C; rom['hE1D]=8'h20; rom['hE1E]=8'h4D; rom['hE1F]=8'h43;
    rom['hE20]=8'h53; rom['hE21]=8'h2D; rom['hE22]=8'h34; rom['hE23]=8'h20;
    rom['hE24]=8'h28; rom['hE25]=8'h34; rom['hE26]=8'h30; rom['hE27]=8'h30;
    rom['hE28]=8'h34; rom['hE29]=8'h29; rom['hE2A]=8'h0D; rom['hE2B]=8'h0A;
    rom['hE2C]=8'h54; rom['hE2D]=8'h69; rom['hE2E]=8'h6E; rom['hE2F]=8'h79;
    rom['hE30]=8'h20; rom['hE31]=8'h4D; rom['hE32]=8'h6F; rom['hE33]=8'h6E;
    rom['hE34]=8'h69; rom['hE35]=8'h74; rom['hE36]=8'h6F; rom['hE37]=8'h72;
    rom['hE38]=8'h0D; rom['hE39]=8'h0A; rom['hE3A]=8'h00; rom['hE3B]=8'h1B;
    rom['hE3C]=8'h40; rom['hE3D]=8'h1F; rom['hE3E]=8'h02; rom['hE3F]=8'h00;
    rom['hE40]=8'h20; rom['hE41]=8'h42; rom['hE42]=8'h41; rom['hE43]=8'h4E;
    rom['hE44]=8'h4B; rom['hE45]=8'h3D; rom['hE46]=8'h00; rom['hE47]=8'h20;
    rom['hE48]=8'h43; rom['hE49]=8'h48; rom['hE4A]=8'h49; rom['hE4B]=8'h50;
    rom['hE4C]=8'h3D; rom['hE4D]=8'h00; rom['hE4E]=8'h20; rom['hE4F]=8'h41;
    rom['hE50]=8'h44; rom['hE51]=8'h52; rom['hE52]=8'h3D; rom['hE53]=8'h00;
    rom['hE54]=8'h0D; rom['hE55]=8'h0A; rom['hE56]=8'h56; rom['hE57]=8'h54;
    rom['hE58]=8'h4C; rom['hE59]=8'h2D; rom['hE5A]=8'h34; rom['hE5B]=8'h30;
    rom['hE5C]=8'h30; rom['hE5D]=8'h34; rom['hE5E]=8'h20; rom['hE5F]=8'h49;
    rom['hE60]=8'h6E; rom['hE61]=8'h74; rom['hE62]=8'h65; rom['hE63]=8'h72;
    rom['hE64]=8'h70; rom['hE65]=8'h72; rom['hE66]=8'h65; rom['hE67]=8'h74;
    rom['hE68]=8'h65; rom['hE69]=8'h72; rom['hE6A]=8'h20; rom['hE6B]=8'h56;
    rom['hE6C]=8'h65; rom['hE6D]=8'h72; rom['hE6E]=8'h20; rom['hE6F]=8'h31;
    rom['hE70]=8'h2E; rom['hE71]=8'h30; rom['hE72]=8'h0D; rom['hE73]=8'h0A;
    rom['hE74]=8'h00; rom['hE75]=8'h0D; rom['hE76]=8'h0A; rom['hE77]=8'h4F;
    rom['hE78]=8'h4B; rom['hE79]=8'h0D; rom['hE7A]=8'h0A; rom['hE7B]=8'h00;
    rom['hE7C]=8'h45; rom['hE7D]=8'h52; rom['hE7E]=8'h52; rom['hE7F]=8'h4F;
    rom['hE80]=8'h52; rom['hE81]=8'h3D; rom['hE82]=8'h00; rom['hE83]=8'h42;
    rom['hE84]=8'h55; rom['hE85]=8'h46; rom['hE86]=8'h3D; rom['hE87]=8'h00;
    rom['hE88]=8'h53; rom['hE89]=8'h50; rom['hE8A]=8'h3D; rom['hE8B]=8'h00;
    rom['hE8C]=8'h49; rom['hE8D]=8'h4E; rom['hE8E]=8'h20; rom['hE8F]=8'h23;
    rom['hE90]=8'h00; rom['hE91]=8'h0D; rom['hE92]=8'h0A; rom['hE93]=8'h76;
    rom['hE94]=8'h3D; rom['hE95]=8'h56; rom['hE96]=8'h54; rom['hE97]=8'h4C;
    rom['hE98]=8'h2C; rom['hE99]=8'h20; rom['hE9A]=8'h72; rom['hE9B]=8'h2F;
    rom['hE9C]=8'h77; rom['hE9D]=8'h3D; rom['hE9E]=8'h52; rom['hE9F]=8'h44;
    rom['hEA0]=8'h2F; rom['hEA1]=8'h57; rom['hEA2]=8'h52; rom['hEA3]=8'h20;
    rom['hEA4]=8'h52; rom['hEA5]=8'h41; rom['hEA6]=8'h4D; rom['hEA7]=8'h2C;
    rom['hEA8]=8'h20; rom['hEA9]=8'h52; rom['hEAA]=8'h2F; rom['hEAB]=8'h57;
    rom['hEAC]=8'h2F; rom['hEAD]=8'h43; rom['hEAE]=8'h2F; rom['hEAF]=8'h42;
    rom['hEB0]=8'h3D; rom['hEB1]=8'h52; rom['hEB2]=8'h44; rom['hEB3]=8'h2F;
    rom['hEB4]=8'h57; rom['hEB5]=8'h52; rom['hEB6]=8'h2F; rom['hEB7]=8'h43;
    rom['hEB8]=8'h4C; rom['hEB9]=8'h52; rom['hEBA]=8'h2F; rom['hEBB]=8'h42;
    rom['hEBC]=8'h4E; rom['hEBD]=8'h4B; rom['hEBE]=8'h20; rom['hEBF]=8'h50;
    rom['hEC0]=8'h4D; rom['hEC1]=8'h2C; rom['hEC2]=8'h20; rom['hEC3]=8'h6C;
    rom['hEC4]=8'h2F; rom['hEC5]=8'h4C; rom['hEC6]=8'h3D; rom['hEC7]=8'h72;
    rom['hEC8]=8'h64; rom['hEC9]=8'h2F; rom['hECA]=8'h77; rom['hECB]=8'h72;
    rom['hECC]=8'h20; rom['hECD]=8'h4C; rom['hECE]=8'h4D; rom['hECF]=8'h2C;
    rom['hED0]=8'h20; rom['hED1]=8'h67; rom['hED2]=8'h3D; rom['hED3]=8'h67;
    rom['hED4]=8'h6F; rom['hED5]=8'h20; rom['hED6]=8'h50; rom['hED7]=8'h4D;
    rom['hED8]=8'h28; rom['hED9]=8'h46; rom['hEDA]=8'h30; rom['hEDB]=8'h30;
    rom['hEDC]=8'h29; rom['hEDD]=8'h0D; rom['hEDE]=8'h0A; rom['hEDF]=8'h00;
    rom['hEE0]=8'h32; rom['hEE1]=8'hC0; rom['hEE2]=8'h00; rom['hEE3]=8'h00;
    rom['hEE4]=8'h00; rom['hEE5]=8'h00; rom['hEE6]=8'h00; rom['hEE7]=8'h00;
    rom['hEE8]=8'h00; rom['hEE9]=8'h00; rom['hEEA]=8'h00; rom['hEEB]=8'h00;
    rom['hEEC]=8'h00; rom['hEED]=8'h00; rom['hEEE]=8'h00; rom['hEEF]=8'h00;
    rom['hEF0]=8'h00; rom['hEF1]=8'h00; rom['hEF2]=8'h00; rom['hEF3]=8'h00;
    rom['hEF4]=8'h00; rom['hEF5]=8'h00; rom['hEF6]=8'h00; rom['hEF7]=8'h00;
    rom['hEF8]=8'h00; rom['hEF9]=8'h00; rom['hEFA]=8'h00; rom['hEFB]=8'h00;
    rom['hEFC]=8'h00; rom['hEFD]=8'h00; rom['hEFE]=8'h00; rom['hEFF]=8'h00;
    rom['hF00]=8'h00; rom['hF01]=8'h00; rom['hF02]=8'h00; rom['hF03]=8'h00;
    rom['hF04]=8'h00; rom['hF05]=8'h00; rom['hF06]=8'h00; rom['hF07]=8'h00;
    rom['hF08]=8'h00; rom['hF09]=8'h00; rom['hF0A]=8'h00; rom['hF0B]=8'h00;
    rom['hF0C]=8'h00; rom['hF0D]=8'h00; rom['hF0E]=8'h00; rom['hF0F]=8'h00;
    rom['hF10]=8'h00; rom['hF11]=8'h00; rom['hF12]=8'h00; rom['hF13]=8'h00;
    rom['hF14]=8'h00; rom['hF15]=8'h00; rom['hF16]=8'h00; rom['hF17]=8'h00;
    rom['hF18]=8'h00; rom['hF19]=8'h00; rom['hF1A]=8'h00; rom['hF1B]=8'h00;
    rom['hF1C]=8'h00; rom['hF1D]=8'h00; rom['hF1E]=8'h00; rom['hF1F]=8'h00;
    rom['hF20]=8'h00; rom['hF21]=8'h00; rom['hF22]=8'h00; rom['hF23]=8'h00;
    rom['hF24]=8'h00; rom['hF25]=8'h00; rom['hF26]=8'h00; rom['hF27]=8'h00;
    rom['hF28]=8'h00; rom['hF29]=8'h00; rom['hF2A]=8'h00; rom['hF2B]=8'h00;
    rom['hF2C]=8'h00; rom['hF2D]=8'h00; rom['hF2E]=8'h00; rom['hF2F]=8'h00;
    rom['hF30]=8'h00; rom['hF31]=8'h00; rom['hF32]=8'h00; rom['hF33]=8'h00;
    rom['hF34]=8'h00; rom['hF35]=8'h00; rom['hF36]=8'h00; rom['hF37]=8'h00;
    rom['hF38]=8'h00; rom['hF39]=8'h00; rom['hF3A]=8'h00; rom['hF3B]=8'h00;
    rom['hF3C]=8'h00; rom['hF3D]=8'h00; rom['hF3E]=8'h00; rom['hF3F]=8'h00;
    rom['hF40]=8'h00; rom['hF41]=8'h00; rom['hF42]=8'h00; rom['hF43]=8'h00;
    rom['hF44]=8'h00; rom['hF45]=8'h00; rom['hF46]=8'h00; rom['hF47]=8'h00;
    rom['hF48]=8'h00; rom['hF49]=8'h00; rom['hF4A]=8'h00; rom['hF4B]=8'h00;
    rom['hF4C]=8'h00; rom['hF4D]=8'h00; rom['hF4E]=8'h00; rom['hF4F]=8'h00;
    rom['hF50]=8'h00; rom['hF51]=8'h00; rom['hF52]=8'h00; rom['hF53]=8'h00;
    rom['hF54]=8'h00; rom['hF55]=8'h00; rom['hF56]=8'h00; rom['hF57]=8'h00;
    rom['hF58]=8'h00; rom['hF59]=8'h00; rom['hF5A]=8'h00; rom['hF5B]=8'h00;
    rom['hF5C]=8'h00; rom['hF5D]=8'h00; rom['hF5E]=8'h00; rom['hF5F]=8'h00;
    rom['hF60]=8'h00; rom['hF61]=8'h00; rom['hF62]=8'h00; rom['hF63]=8'h00;
    rom['hF64]=8'h00; rom['hF65]=8'h00; rom['hF66]=8'h00; rom['hF67]=8'h00;
    rom['hF68]=8'h00; rom['hF69]=8'h00; rom['hF6A]=8'h00; rom['hF6B]=8'h00;
    rom['hF6C]=8'h00; rom['hF6D]=8'h00; rom['hF6E]=8'h00; rom['hF6F]=8'h00;
    rom['hF70]=8'h00; rom['hF71]=8'h00; rom['hF72]=8'h00; rom['hF73]=8'h00;
    rom['hF74]=8'h00; rom['hF75]=8'h00; rom['hF76]=8'h00; rom['hF77]=8'h00;
    rom['hF78]=8'h00; rom['hF79]=8'h00; rom['hF7A]=8'h00; rom['hF7B]=8'h00;
    rom['hF7C]=8'h00; rom['hF7D]=8'h00; rom['hF7E]=8'h00; rom['hF7F]=8'h00;
    rom['hF80]=8'h00; rom['hF81]=8'h00; rom['hF82]=8'h00; rom['hF83]=8'h00;
    rom['hF84]=8'h00; rom['hF85]=8'h00; rom['hF86]=8'h00; rom['hF87]=8'h00;
    rom['hF88]=8'h00; rom['hF89]=8'h00; rom['hF8A]=8'h00; rom['hF8B]=8'h00;
    rom['hF8C]=8'h00; rom['hF8D]=8'h00; rom['hF8E]=8'h00; rom['hF8F]=8'h00;
    rom['hF90]=8'h00; rom['hF91]=8'h00; rom['hF92]=8'h00; rom['hF93]=8'h00;
    rom['hF94]=8'h00; rom['hF95]=8'h00; rom['hF96]=8'h00; rom['hF97]=8'h00;
    rom['hF98]=8'h00; rom['hF99]=8'h00; rom['hF9A]=8'h00; rom['hF9B]=8'h00;
    rom['hF9C]=8'h00; rom['hF9D]=8'h00; rom['hF9E]=8'h00; rom['hF9F]=8'h00;
    rom['hFA0]=8'h00; rom['hFA1]=8'h00; rom['hFA2]=8'h00; rom['hFA3]=8'h00;
    rom['hFA4]=8'h00; rom['hFA5]=8'h00; rom['hFA6]=8'h00; rom['hFA7]=8'h00;
    rom['hFA8]=8'h00; rom['hFA9]=8'h00; rom['hFAA]=8'h00; rom['hFAB]=8'h00;
    rom['hFAC]=8'h00; rom['hFAD]=8'h00; rom['hFAE]=8'h00; rom['hFAF]=8'h00;
    rom['hFB0]=8'h00; rom['hFB1]=8'h00; rom['hFB2]=8'h00; rom['hFB3]=8'h00;
    rom['hFB4]=8'h00; rom['hFB5]=8'h00; rom['hFB6]=8'h00; rom['hFB7]=8'h00;
    rom['hFB8]=8'h00; rom['hFB9]=8'h00; rom['hFBA]=8'h00; rom['hFBB]=8'h00;
    rom['hFBC]=8'h00; rom['hFBD]=8'h00; rom['hFBE]=8'h00; rom['hFBF]=8'h00;
    rom['hFC0]=8'h00; rom['hFC1]=8'h00; rom['hFC2]=8'h00; rom['hFC3]=8'h00;
    rom['hFC4]=8'h00; rom['hFC5]=8'h00; rom['hFC6]=8'h00; rom['hFC7]=8'h00;
    rom['hFC8]=8'h00; rom['hFC9]=8'h00; rom['hFCA]=8'h00; rom['hFCB]=8'h00;
    rom['hFCC]=8'h00; rom['hFCD]=8'h00; rom['hFCE]=8'h00; rom['hFCF]=8'h00;
    rom['hFD0]=8'h00; rom['hFD1]=8'h00; rom['hFD2]=8'h00; rom['hFD3]=8'h00;
    rom['hFD4]=8'h00; rom['hFD5]=8'h00; rom['hFD6]=8'h00; rom['hFD7]=8'h00;
    rom['hFD8]=8'h00; rom['hFD9]=8'h00; rom['hFDA]=8'h00; rom['hFDB]=8'h00;
    rom['hFDC]=8'h00; rom['hFDD]=8'h00; rom['hFDE]=8'h00; rom['hFDF]=8'h00;
    rom['hFE0]=8'h00; rom['hFE1]=8'h00; rom['hFE2]=8'h00; rom['hFE3]=8'h00;
    rom['hFE4]=8'h00; rom['hFE5]=8'h00; rom['hFE6]=8'h00; rom['hFE7]=8'h00;
    rom['hFE8]=8'h00; rom['hFE9]=8'h00; rom['hFEA]=8'h00; rom['hFEB]=8'h00;
    rom['hFEC]=8'h00; rom['hFED]=8'h00; rom['hFEE]=8'h00; rom['hFEF]=8'h00;
    rom['hFF0]=8'h00; rom['hFF1]=8'h00; rom['hFF2]=8'h00; rom['hFF3]=8'h00;
    rom['hFF4]=8'h00; rom['hFF5]=8'h00; rom['hFF6]=8'h00; rom['hFF7]=8'h00;
    rom['hFF8]=8'h00; rom['hFF9]=8'h00; rom['hFFA]=8'h00; rom['hFFB]=8'h00;
    rom['hFFC]=8'h00; rom['hFFD]=8'h00; rom['hFFE]=8'h00; rom['hFFF]=8'h00;

    end
endmodule
