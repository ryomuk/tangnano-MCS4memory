//-----------------------------------------------------------------------------
//
// ROM image
//
//-----------------------------------------------------------------------------
module rom_image( addr, dout );
//-----------------------------------------------------------------------------
  input [11:0] addr;
  output [7:0] dout;
//-----------------------------------------------------------------------------
  reg [7:0]    rom [4095:0];
//-----------------------------------------------------------------------------
  assign dout = rom[addr];
  initial
    begin
       //
       // place rom data here
       //
    end
endmodule
