//-----------------------------------------------------------------------------
//
// ROM image
//
//-----------------------------------------------------------------------------
module rom_image( addr, dout );
//-----------------------------------------------------------------------------
  input [11:0] addr;
  output [7:0] dout;
//-----------------------------------------------------------------------------
  reg [7:0]    rom [4095:0];
//-----------------------------------------------------------------------------
  assign dout = rom[addr];
  initial
    begin
    rom['h000]=8'h00; rom['h001]=8'hF0; rom['h002]=8'hFD; rom['h003]=8'h28;
    rom['h004]=8'h80; rom['h005]=8'h5C; rom['h006]=8'h7F; rom['h007]=8'hD0;
    rom['h008]=8'hB2; rom['h009]=8'hD0; rom['h00A]=8'hB3; rom['h00B]=8'h5B;
    rom['h00C]=8'hB9; rom['h00D]=8'h5B; rom['h00E]=8'hAD; rom['h00F]=8'h73;
    rom['h010]=8'h0B; rom['h011]=8'h72; rom['h012]=8'h09; rom['h013]=8'h22;
    rom['h014]=8'h00; rom['h015]=8'h5B; rom['h016]=8'hB9; rom['h017]=8'h20;
    rom['h018]=8'h42; rom['h019]=8'h5E; rom['h01A]=8'h00; rom['h01B]=8'h20;
    rom['h01C]=8'h1F; rom['h01D]=8'h5E; rom['h01E]=8'h00; rom['h01F]=8'h20;
    rom['h020]=8'h38; rom['h021]=8'h22; rom['h022]=8'h44; rom['h023]=8'h57;
    rom['h024]=8'hF1; rom['h025]=8'h20; rom['h026]=8'h14; rom['h027]=8'h24;
    rom['h028]=8'h00; rom['h029]=8'h26; rom['h02A]=8'h00; rom['h02B]=8'h57;
    rom['h02C]=8'h96; rom['h02D]=8'h22; rom['h02E]=8'h5D; rom['h02F]=8'h5C;
    rom['h030]=8'h5F; rom['h031]=8'h20; rom['h032]=8'h28; rom['h033]=8'h24;
    rom['h034]=8'hFD; rom['h035]=8'h26; rom['h036]=8'h00; rom['h037]=8'h57;
    rom['h038]=8'h96; rom['h039]=8'h5B; rom['h03A]=8'hC4; rom['h03B]=8'h5B;
    rom['h03C]=8'h5D; rom['h03D]=8'h5D; rom['h03E]=8'h4B; rom['h03F]=8'h2E;
    rom['h040]=8'h48; rom['h041]=8'h5D; rom['h042]=8'h27; rom['h043]=8'h1C;
    rom['h044]=8'h47; rom['h045]=8'h40; rom['h046]=8'hE9; rom['h047]=8'h2E;
    rom['h048]=8'h44; rom['h049]=8'h5D; rom['h04A]=8'h27; rom['h04B]=8'h1C;
    rom['h04C]=8'h4F; rom['h04D]=8'h40; rom['h04E]=8'h92; rom['h04F]=8'h2E;
    rom['h050]=8'h4C; rom['h051]=8'h5D; rom['h052]=8'h27; rom['h053]=8'h1C;
    rom['h054]=8'h57; rom['h055]=8'h41; rom['h056]=8'h09; rom['h057]=8'h2E;
    rom['h058]=8'h43; rom['h059]=8'h5D; rom['h05A]=8'h27; rom['h05B]=8'h1C;
    rom['h05C]=8'h5F; rom['h05D]=8'h41; rom['h05E]=8'h7B; rom['h05F]=8'h2E;
    rom['h060]=8'h47; rom['h061]=8'h5D; rom['h062]=8'h27; rom['h063]=8'h1C;
    rom['h064]=8'h67; rom['h065]=8'h40; rom['h066]=8'hE7; rom['h067]=8'h2E;
    rom['h068]=8'h45; rom['h069]=8'h5D; rom['h06A]=8'h27; rom['h06B]=8'h1C;
    rom['h06C]=8'h8C; rom['h06D]=8'h5B; rom['h06E]=8'h5D; rom['h06F]=8'h5D;
    rom['h070]=8'h4B; rom['h071]=8'h2E; rom['h072]=8'h53; rom['h073]=8'h5D;
    rom['h074]=8'h27; rom['h075]=8'h1C; rom['h076]=8'h7A; rom['h077]=8'hD2;
    rom['h078]=8'h40; rom['h079]=8'h86; rom['h07A]=8'h2E; rom['h07B]=8'h56;
    rom['h07C]=8'h5D; rom['h07D]=8'h27; rom['h07E]=8'h1C; rom['h07F]=8'h83;
    rom['h080]=8'hD1; rom['h081]=8'h40; rom['h082]=8'h86; rom['h083]=8'h58;
    rom['h084]=8'h6B; rom['h085]=8'hD0; rom['h086]=8'h2E; rom['h087]=8'h24;
    rom['h088]=8'h2F; rom['h089]=8'hE0; rom['h08A]=8'h41; rom['h08B]=8'h95;
    rom['h08C]=8'h20; rom['h08D]=8'h47; rom['h08E]=8'h5E; rom['h08F]=8'h00;
    rom['h090]=8'h40; rom['h091]=8'h2D; rom['h092]=8'h22; rom['h093]=8'h2C;
    rom['h094]=8'h58; rom['h095]=8'hC9; rom['h096]=8'h2E; rom['h097]=8'h38;
    rom['h098]=8'h58; rom['h099]=8'h09; rom['h09A]=8'h2E; rom['h09B]=8'h44;
    rom['h09C]=8'h5D; rom['h09D]=8'h27; rom['h09E]=8'h1C; rom['h09F]=8'hA2;
    rom['h0A0]=8'h40; rom['h0A1]=8'hCE; rom['h0A2]=8'h2E; rom['h0A3]=8'h4C;
    rom['h0A4]=8'h5D; rom['h0A5]=8'h27; rom['h0A6]=8'h1C; rom['h0A7]=8'hAA;
    rom['h0A8]=8'h40; rom['h0A9]=8'hB0; rom['h0AA]=8'h20; rom['h0AB]=8'h4B;
    rom['h0AC]=8'h5E; rom['h0AD]=8'h00; rom['h0AE]=8'h40; rom['h0AF]=8'h2D;
    rom['h0B0]=8'h20; rom['h0B1]=8'h2C; rom['h0B2]=8'h58; rom['h0B3]=8'h11;
    rom['h0B4]=8'hA2; rom['h0B5]=8'hBA; rom['h0B6]=8'hA3; rom['h0B7]=8'hBB;
    rom['h0B8]=8'hD8; rom['h0B9]=8'hBA; rom['h0BA]=8'h22; rom['h0BB]=8'h2C;
    rom['h0BC]=8'h58; rom['h0BD]=8'h29; rom['h0BE]=8'h22; rom['h0BF]=8'h3A;
    rom['h0C0]=8'h5C; rom['h0C1]=8'h5F; rom['h0C2]=8'h5B; rom['h0C3]=8'h5D;
    rom['h0C4]=8'h5C; rom['h0C5]=8'h85; rom['h0C6]=8'h7B; rom['h0C7]=8'hC2;
    rom['h0C8]=8'h5C; rom['h0C9]=8'hA0; rom['h0CA]=8'h7A; rom['h0CB]=8'hBA;
    rom['h0CC]=8'h40; rom['h0CD]=8'h2D; rom['h0CE]=8'h2E; rom['h0CF]=8'h2C;
    rom['h0D0]=8'h58; rom['h0D1]=8'h09; rom['h0D2]=8'hA2; rom['h0D3]=8'hB0;
    rom['h0D4]=8'hA3; rom['h0D5]=8'hB1; rom['h0D6]=8'hDC; rom['h0D7]=8'hBA;
    rom['h0D8]=8'h5D; rom['h0D9]=8'h57; rom['h0DA]=8'h60; rom['h0DB]=8'h7A;
    rom['h0DC]=8'hD8; rom['h0DD]=8'hA0; rom['h0DE]=8'hB2; rom['h0DF]=8'hA1;
    rom['h0E0]=8'hB3; rom['h0E1]=8'h20; rom['h0E2]=8'h2C; rom['h0E3]=8'h57;
    rom['h0E4]=8'hF1; rom['h0E5]=8'h40; rom['h0E6]=8'h2D; rom['h0E7]=8'h4F;
    rom['h0E8]=8'h00; rom['h0E9]=8'h5B; rom['h0EA]=8'h5D; rom['h0EB]=8'h5D;
    rom['h0EC]=8'h34; rom['h0ED]=8'h1C; rom['h0EE]=8'hF1; rom['h0EF]=8'h40;
    rom['h0F0]=8'hFB; rom['h0F1]=8'h5D; rom['h0F2]=8'h4B; rom['h0F3]=8'h24;
    rom['h0F4]=8'h38; rom['h0F5]=8'h57; rom['h0F6]=8'hFD; rom['h0F7]=8'h22;
    rom['h0F8]=8'h2C; rom['h0F9]=8'h58; rom['h0FA]=8'hC9; rom['h0FB]=8'h2E;
    rom['h0FC]=8'h38; rom['h0FD]=8'h58; rom['h0FE]=8'h09; rom['h0FF]=8'h5C;
    rom['h100]=8'h5F; rom['h101]=8'h22; rom['h102]=8'h2C; rom['h103]=8'h58;
    rom['h104]=8'h29; rom['h105]=8'h5C; rom['h106]=8'hA0; rom['h107]=8'h40;
    rom['h108]=8'h2D; rom['h109]=8'h20; rom['h10A]=8'h28; rom['h10B]=8'h24;
    rom['h10C]=8'hFD; rom['h10D]=8'h26; rom['h10E]=8'h00; rom['h10F]=8'h57;
    rom['h110]=8'h96; rom['h111]=8'h5B; rom['h112]=8'hC4; rom['h113]=8'h5B;
    rom['h114]=8'h5D; rom['h115]=8'h5D; rom['h116]=8'h34; rom['h117]=8'h1C;
    rom['h118]=8'h1B; rom['h119]=8'h41; rom['h11A]=8'h73; rom['h11B]=8'h2E;
    rom['h11C]=8'h3A; rom['h11D]=8'h5D; rom['h11E]=8'h27; rom['h11F]=8'h14;
    rom['h120]=8'h23; rom['h121]=8'h41; rom['h122]=8'h49; rom['h123]=8'h5C;
    rom['h124]=8'h18; rom['h125]=8'hA2; rom['h126]=8'hBA; rom['h127]=8'hA3;
    rom['h128]=8'hBB; rom['h129]=8'h5C; rom['h12A]=8'h18; rom['h12B]=8'hA2;
    rom['h12C]=8'hB4; rom['h12D]=8'hA3; rom['h12E]=8'hB5; rom['h12F]=8'h5C;
    rom['h130]=8'h18; rom['h131]=8'hA2; rom['h132]=8'hB6; rom['h133]=8'hA3;
    rom['h134]=8'hB7; rom['h135]=8'h22; rom['h136]=8'h2C; rom['h137]=8'h57;
    rom['h138]=8'h90; rom['h139]=8'h5C; rom['h13A]=8'h18; rom['h13B]=8'h5D;
    rom['h13C]=8'h34; rom['h13D]=8'h1C; rom['h13E]=8'h41; rom['h13F]=8'h41;
    rom['h140]=8'h53; rom['h141]=8'h2E; rom['h142]=8'h01; rom['h143]=8'h5D;
    rom['h144]=8'h27; rom['h145]=8'h1C; rom['h146]=8'h49; rom['h147]=8'h41;
    rom['h148]=8'h73; rom['h149]=8'h58; rom['h14A]=8'h6B; rom['h14B]=8'h5C;
    rom['h14C]=8'h0A; rom['h14D]=8'h20; rom['h14E]=8'h57; rom['h14F]=8'h5E;
    rom['h150]=8'h00; rom['h151]=8'h40; rom['h152]=8'h2D; rom['h153]=8'hAB;
    rom['h154]=8'h1C; rom['h155]=8'h5B; rom['h156]=8'hAA; rom['h157]=8'h1C;
    rom['h158]=8'h5B; rom['h159]=8'h41; rom['h15A]=8'h09; rom['h15B]=8'h20;
    rom['h15C]=8'h28; rom['h15D]=8'h5C; rom['h15E]=8'h18; rom['h15F]=8'h14;
    rom['h160]=8'h63; rom['h161]=8'h41; rom['h162]=8'h09; rom['h163]=8'h20;
    rom['h164]=8'h2C; rom['h165]=8'h5B; rom['h166]=8'h81; rom['h167]=8'h58;
    rom['h168]=8'h5B; rom['h169]=8'hAB; rom['h16A]=8'hF8; rom['h16B]=8'hBB;
    rom['h16C]=8'h12; rom['h16D]=8'h71; rom['h16E]=8'hAA; rom['h16F]=8'hF8;
    rom['h170]=8'hBA; rom['h171]=8'h41; rom['h172]=8'h53; rom['h173]=8'h20;
    rom['h174]=8'h38; rom['h175]=8'h22; rom['h176]=8'h4C; rom['h177]=8'h57;
    rom['h178]=8'hF1; rom['h179]=8'h40; rom['h17A]=8'h2D; rom['h17B]=8'h2A;
    rom['h17C]=8'h00; rom['h17D]=8'hAA; rom['h17E]=8'hB2; rom['h17F]=8'hAB;
    rom['h180]=8'hB3; rom['h181]=8'h5B; rom['h182]=8'hB9; rom['h183]=8'h20;
    rom['h184]=8'h00; rom['h185]=8'h22; rom['h186]=8'h00; rom['h187]=8'h5B;
    rom['h188]=8'hA1; rom['h189]=8'h71; rom['h18A]=8'h87; rom['h18B]=8'h70;
    rom['h18C]=8'h87; rom['h18D]=8'h5B; rom['h18E]=8'hAD; rom['h18F]=8'h7B;
    rom['h190]=8'h7D; rom['h191]=8'h7A; rom['h192]=8'h7D; rom['h193]=8'h40;
    rom['h194]=8'h2D; rom['h195]=8'h22; rom['h196]=8'h14; rom['h197]=8'h58;
    rom['h198]=8'hC9; rom['h199]=8'h20; rom['h19A]=8'h65; rom['h19B]=8'h5E;
    rom['h19C]=8'h00; rom['h19D]=8'h2E; rom['h19E]=8'h24; rom['h19F]=8'h2F;
    rom['h1A0]=8'hE9; rom['h1A1]=8'h14; rom['h1A2]=8'hA5; rom['h1A3]=8'h41;
    rom['h1A4]=8'hBB; rom['h1A5]=8'h51; rom['h1A6]=8'hE6; rom['h1A7]=8'h11;
    rom['h1A8]=8'hAB; rom['h1A9]=8'h41; rom['h1AA]=8'hA5; rom['h1AB]=8'h2A;
    rom['h1AC]=8'h00; rom['h1AD]=8'h19; rom['h1AE]=8'hA5; rom['h1AF]=8'h7B;
    rom['h1B0]=8'hAD; rom['h1B1]=8'h7A; rom['h1B2]=8'hAD; rom['h1B3]=8'h11;
    rom['h1B4]=8'hB3; rom['h1B5]=8'h20; rom['h1B6]=8'hC2; rom['h1B7]=8'h5E;
    rom['h1B8]=8'h00; rom['h1B9]=8'h42; rom['h1BA]=8'h6B; rom['h1BB]=8'hF8;
    rom['h1BC]=8'h14; rom['h1BD]=8'hC0; rom['h1BE]=8'h41; rom['h1BF]=8'hD4;
    rom['h1C0]=8'h20; rom['h1C1]=8'h87; rom['h1C2]=8'h5E; rom['h1C3]=8'h00;
    rom['h1C4]=8'h5C; rom['h1C5]=8'hAC; rom['h1C6]=8'h58; rom['h1C7]=8'hEE;
    rom['h1C8]=8'h11; rom['h1C9]=8'hCE; rom['h1CA]=8'h51; rom['h1CB]=8'hE6;
    rom['h1CC]=8'h41; rom['h1CD]=8'hC4; rom['h1CE]=8'h11; rom['h1CF]=8'hCE;
    rom['h1D0]=8'h5C; rom['h1D1]=8'hA0; rom['h1D2]=8'h40; rom['h1D3]=8'h2D;
    rom['h1D4]=8'h58; rom['h1D5]=8'hEA; rom['h1D6]=8'h5C; rom['h1D7]=8'hA0;
    rom['h1D8]=8'h5C; rom['h1D9]=8'h37; rom['h1DA]=8'h2E; rom['h1DB]=8'h2E;
    rom['h1DC]=8'h5D; rom['h1DD]=8'h27; rom['h1DE]=8'h14; rom['h1DF]=8'hE4;
    rom['h1E0]=8'h51; rom['h1E1]=8'hE6; rom['h1E2]=8'h41; rom['h1E3]=8'hD4;
    rom['h1E4]=8'h40; rom['h1E5]=8'h2D; rom['h1E6]=8'h20; rom['h1E7]=8'h14;
    rom['h1E8]=8'h5B; rom['h1E9]=8'h5D; rom['h1EA]=8'hA2; rom['h1EB]=8'hF5;
    rom['h1EC]=8'h1A; rom['h1ED]=8'hF0; rom['h1EE]=8'h42; rom['h1EF]=8'h06;
    rom['h1F0]=8'hF5; rom['h1F1]=8'h1A; rom['h1F2]=8'hF5; rom['h1F3]=8'h42;
    rom['h1F4]=8'h0B; rom['h1F5]=8'hA3; rom['h1F6]=8'h1C; rom['h1F7]=8'hFD;
    rom['h1F8]=8'hA2; rom['h1F9]=8'h1C; rom['h1FA]=8'hFD; rom['h1FB]=8'h42;
    rom['h1FC]=8'h71; rom['h1FD]=8'hA3; rom['h1FE]=8'hF1; rom['h1FF]=8'hF5;
    rom['h200]=8'hB3; rom['h201]=8'hA2; rom['h202]=8'hF5; rom['h203]=8'hB2;
    rom['h204]=8'h4A; rom['h205]=8'h00; rom['h206]=8'hF5; rom['h207]=8'h1A;
    rom['h208]=8'h0B; rom['h209]=8'h41; rom['h20A]=8'hFD; rom['h20B]=8'h5B;
    rom['h20C]=8'h12; rom['h20D]=8'hF0; rom['h20E]=8'hB2; rom['h20F]=8'hA3;
    rom['h210]=8'hF4; rom['h211]=8'hF1; rom['h212]=8'hF5; rom['h213]=8'hB3;
    rom['h214]=8'hA3; rom['h215]=8'hD2; rom['h216]=8'hF1; rom['h217]=8'h93;
    rom['h218]=8'h14; rom['h219]=8'h1E; rom['h21A]=8'h58; rom['h21B]=8'h17;
    rom['h21C]=8'h42; rom['h21D]=8'h24; rom['h21E]=8'h20; rom['h21F]=8'h04;
    rom['h220]=8'h5B; rom['h221]=8'h5D; rom['h222]=8'h58; rom['h223]=8'h6B;
    rom['h224]=8'h20; rom['h225]=8'h12; rom['h226]=8'h57; rom['h227]=8'hF1;
    rom['h228]=8'h5B; rom['h229]=8'h43; rom['h22A]=8'hA2; rom['h22B]=8'hF5;
    rom['h22C]=8'h1A; rom['h22D]=8'h30; rom['h22E]=8'h42; rom['h22F]=8'h58;
    rom['h230]=8'h2E; rom['h231]=8'h76; rom['h232]=8'h5D; rom['h233]=8'h27;
    rom['h234]=8'h1C; rom['h235]=8'h38; rom['h236]=8'h42; rom['h237]=8'h67;
    rom['h238]=8'h24; rom['h239]=8'h00; rom['h23A]=8'hA2; rom['h23B]=8'hF5;
    rom['h23C]=8'hF5; rom['h23D]=8'hF1; rom['h23E]=8'hF6; rom['h23F]=8'hF6;
    rom['h240]=8'hB5; rom['h241]=8'hA3; rom['h242]=8'hF5; rom['h243]=8'hA5;
    rom['h244]=8'hF5; rom['h245]=8'hF4; rom['h246]=8'hF5; rom['h247]=8'hB5;
    rom['h248]=8'h22; rom['h249]=8'h12; rom['h24A]=8'h58; rom['h24B]=8'h17;
    rom['h24C]=8'hD2; rom['h24D]=8'hF1; rom['h24E]=8'h95; rom['h24F]=8'h14;
    rom['h250]=8'h54; rom['h251]=8'h57; rom['h252]=8'hFD; rom['h253]=8'hC0;
    rom['h254]=8'h20; rom['h255]=8'h04; rom['h256]=8'h4B; rom['h257]=8'h81;
    rom['h258]=8'h24; rom['h259]=8'hF0; rom['h25A]=8'hA3; rom['h25B]=8'hF5;
    rom['h25C]=8'hA2; rom['h25D]=8'hF5; rom['h25E]=8'hF1; rom['h25F]=8'hF5;
    rom['h260]=8'hB5; rom['h261]=8'h2E; rom['h262]=8'h12; rom['h263]=8'h58;
    rom['h264]=8'h09; rom['h265]=8'h49; rom['h266]=8'hEF; rom['h267]=8'h20;
    rom['h268]=8'hCB; rom['h269]=8'h5E; rom['h26A]=8'h00; rom['h26B]=8'h58;
    rom['h26C]=8'hEA; rom['h26D]=8'h5C; rom['h26E]=8'hA0; rom['h26F]=8'h40;
    rom['h270]=8'h2D; rom['h271]=8'hC0; rom['h272]=8'h5B; rom['h273]=8'h5D;
    rom['h274]=8'h24; rom['h275]=8'h0C; rom['h276]=8'h57; rom['h277]=8'hFD;
    rom['h278]=8'h5B; rom['h279]=8'h5D; rom['h27A]=8'h24; rom['h27B]=8'h0E;
    rom['h27C]=8'h47; rom['h27D]=8'hFD; rom['h27E]=8'h2E; rom['h27F]=8'h00;
    rom['h280]=8'h58; rom['h281]=8'h09; rom['h282]=8'h20; rom['h283]=8'h0C;
    rom['h284]=8'h4B; rom['h285]=8'h81; rom['h286]=8'h20; rom['h287]=8'h0C;
    rom['h288]=8'h48; rom['h289]=8'h5B; rom['h28A]=8'h22; rom['h28B]=8'h0E;
    rom['h28C]=8'h44; rom['h28D]=8'h30; rom['h28E]=8'h22; rom['h28F]=8'h0E;
    rom['h290]=8'h44; rom['h291]=8'h36; rom['h292]=8'h24; rom['h293]=8'h0E;
    rom['h294]=8'h44; rom['h295]=8'h3C; rom['h296]=8'h20; rom['h297]=8'h00;
    rom['h298]=8'h58; rom['h299]=8'h11; rom['h29A]=8'hA2; rom['h29B]=8'hF5;
    rom['h29C]=8'hA3; rom['h29D]=8'hF5; rom['h29E]=8'hB3; rom['h29F]=8'hA2;
    rom['h2A0]=8'hF5; rom['h2A1]=8'hB2; rom['h2A2]=8'h56; rom['h2A3]=8'h8C;
    rom['h2A4]=8'h47; rom['h2A5]=8'hF1; rom['h2A6]=8'hC0; rom['h2A7]=8'h20;
    rom['h2A8]=8'h04; rom['h2A9]=8'h22; rom['h2AA]=8'h0C; rom['h2AB]=8'h58;
    rom['h2AC]=8'hA0; rom['h2AD]=8'h46; rom['h2AE]=8'h8C; rom['h2AF]=8'h20;
    rom['h2B0]=8'h0C; rom['h2B1]=8'h5B; rom['h2B2]=8'h5D; rom['h2B3]=8'h58;
    rom['h2B4]=8'h6B; rom['h2B5]=8'h24; rom['h2B6]=8'h00; rom['h2B7]=8'h47;
    rom['h2B8]=8'hFD; rom['h2B9]=8'h20; rom['h2BA]=8'h0C; rom['h2BB]=8'h48;
    rom['h2BC]=8'h6B; rom['h2BD]=8'h22; rom['h2BE]=8'h0C; rom['h2BF]=8'h44;
    rom['h2C0]=8'h30; rom['h2C1]=8'h22; rom['h2C2]=8'h0C; rom['h2C3]=8'h44;
    rom['h2C4]=8'h36; rom['h2C5]=8'h24; rom['h2C6]=8'h0C; rom['h2C7]=8'h44;
    rom['h2C8]=8'h3C; rom['h2C9]=8'h20; rom['h2CA]=8'h00; rom['h2CB]=8'h58;
    rom['h2CC]=8'h11; rom['h2CD]=8'hA3; rom['h2CE]=8'hF6; rom['h2CF]=8'hA2;
    rom['h2D0]=8'hF6; rom['h2D1]=8'hB2; rom['h2D2]=8'hA3; rom['h2D3]=8'hF6;
    rom['h2D4]=8'hB3; rom['h2D5]=8'h56; rom['h2D6]=8'h8C; rom['h2D7]=8'h47;
    rom['h2D8]=8'hF1; rom['h2D9]=8'hC0; rom['h2DA]=8'h5B; rom['h2DB]=8'h5D;
    rom['h2DC]=8'h24; rom['h2DD]=8'h08; rom['h2DE]=8'h57; rom['h2DF]=8'hFD;
    rom['h2E0]=8'h5B; rom['h2E1]=8'h5D; rom['h2E2]=8'h24; rom['h2E3]=8'h0A;
    rom['h2E4]=8'h47; rom['h2E5]=8'hFD; rom['h2E6]=8'h2E; rom['h2E7]=8'h00;
    rom['h2E8]=8'h58; rom['h2E9]=8'h09; rom['h2EA]=8'h20; rom['h2EB]=8'h08;
    rom['h2EC]=8'h4B; rom['h2ED]=8'h81; rom['h2EE]=8'h20; rom['h2EF]=8'h08;
    rom['h2F0]=8'h48; rom['h2F1]=8'h5B; rom['h2F2]=8'h22; rom['h2F3]=8'h0A;
    rom['h2F4]=8'h44; rom['h2F5]=8'h30; rom['h2F6]=8'h22; rom['h2F7]=8'h0A;
    rom['h2F8]=8'h44; rom['h2F9]=8'h36; rom['h2FA]=8'h24; rom['h2FB]=8'h0A;
    rom['h2FC]=8'h44; rom['h2FD]=8'h3C; rom['h2FE]=8'h20; rom['h2FF]=8'h00;
    rom['h300]=8'h58; rom['h301]=8'h11; rom['h302]=8'h56; rom['h303]=8'h40;
    rom['h304]=8'hA3; rom['h305]=8'hF5; rom['h306]=8'hB3; rom['h307]=8'hA2;
    rom['h308]=8'hF5; rom['h309]=8'hB2; rom['h30A]=8'h56; rom['h30B]=8'h8C;
    rom['h30C]=8'h47; rom['h30D]=8'hF1; rom['h30E]=8'hC0; rom['h30F]=8'h20;
    rom['h310]=8'h04; rom['h311]=8'h22; rom['h312]=8'h08; rom['h313]=8'h58;
    rom['h314]=8'hA0; rom['h315]=8'h46; rom['h316]=8'h8C; rom['h317]=8'h20;
    rom['h318]=8'h08; rom['h319]=8'h5B; rom['h31A]=8'h5D; rom['h31B]=8'h58;
    rom['h31C]=8'h6B; rom['h31D]=8'h24; rom['h31E]=8'h00; rom['h31F]=8'h47;
    rom['h320]=8'hFD; rom['h321]=8'h20; rom['h322]=8'h08; rom['h323]=8'h48;
    rom['h324]=8'h6B; rom['h325]=8'h22; rom['h326]=8'h08; rom['h327]=8'h44;
    rom['h328]=8'h30; rom['h329]=8'h22; rom['h32A]=8'h08; rom['h32B]=8'h44;
    rom['h32C]=8'h36; rom['h32D]=8'h24; rom['h32E]=8'h08; rom['h32F]=8'h44;
    rom['h330]=8'h3C; rom['h331]=8'h20; rom['h332]=8'h00; rom['h333]=8'h58;
    rom['h334]=8'h11; rom['h335]=8'h56; rom['h336]=8'h40; rom['h337]=8'hA2;
    rom['h338]=8'hF6; rom['h339]=8'hB2; rom['h33A]=8'hA3; rom['h33B]=8'hF6;
    rom['h33C]=8'hB3; rom['h33D]=8'h56; rom['h33E]=8'h8C; rom['h33F]=8'h47;
    rom['h340]=8'hF1; rom['h341]=8'hC0; rom['h342]=8'h5B; rom['h343]=8'h5D;
    rom['h344]=8'h24; rom['h345]=8'h04; rom['h346]=8'h57; rom['h347]=8'hFD;
    rom['h348]=8'h5B; rom['h349]=8'h5D; rom['h34A]=8'h24; rom['h34B]=8'h06;
    rom['h34C]=8'h47; rom['h34D]=8'hFD; rom['h34E]=8'h5B; rom['h34F]=8'h5D;
    rom['h350]=8'h24; rom['h351]=8'h1C; rom['h352]=8'h57; rom['h353]=8'hFD;
    rom['h354]=8'h5B; rom['h355]=8'h5D; rom['h356]=8'h24; rom['h357]=8'h1E;
    rom['h358]=8'h57; rom['h359]=8'hFD; rom['h35A]=8'h2E; rom['h35B]=8'h04;
    rom['h35C]=8'h58; rom['h35D]=8'h09; rom['h35E]=8'h20; rom['h35F]=8'h1C;
    rom['h360]=8'h5B; rom['h361]=8'h81; rom['h362]=8'h58; rom['h363]=8'h5B;
    rom['h364]=8'h2E; rom['h365]=8'h06; rom['h366]=8'h58; rom['h367]=8'h09;
    rom['h368]=8'h5B; rom['h369]=8'h81; rom['h36A]=8'h48; rom['h36B]=8'h5B;
    rom['h36C]=8'h20; rom['h36D]=8'h04; rom['h36E]=8'h48; rom['h36F]=8'h5B;
    rom['h370]=8'h22; rom['h371]=8'h06; rom['h372]=8'h44; rom['h373]=8'h30;
    rom['h374]=8'h22; rom['h375]=8'h06; rom['h376]=8'h44; rom['h377]=8'h36;
    rom['h378]=8'h24; rom['h379]=8'h06; rom['h37A]=8'h44; rom['h37B]=8'h3C;
    rom['h37C]=8'h20; rom['h37D]=8'h00; rom['h37E]=8'h58; rom['h37F]=8'h11;
    rom['h380]=8'hA3; rom['h381]=8'hFB; rom['h382]=8'hB3; rom['h383]=8'hD0;
    rom['h384]=8'h82; rom['h385]=8'hFB; rom['h386]=8'hB2; rom['h387]=8'h47;
    rom['h388]=8'hF1; rom['h389]=8'hC0; rom['h38A]=8'h20; rom['h38B]=8'h04;
    rom['h38C]=8'h22; rom['h38D]=8'h04; rom['h38E]=8'h58; rom['h38F]=8'hA0;
    rom['h390]=8'h46; rom['h391]=8'h8C; rom['h392]=8'h5B; rom['h393]=8'h5D;
    rom['h394]=8'h24; rom['h395]=8'h1C; rom['h396]=8'h57; rom['h397]=8'hFD;
    rom['h398]=8'h5B; rom['h399]=8'h5D; rom['h39A]=8'h24; rom['h39B]=8'h1E;
    rom['h39C]=8'h57; rom['h39D]=8'hFD; rom['h39E]=8'h20; rom['h39F]=8'h1C;
    rom['h3A0]=8'h24; rom['h3A1]=8'h04; rom['h3A2]=8'h5B; rom['h3A3]=8'h5D;
    rom['h3A4]=8'h57; rom['h3A5]=8'hFD; rom['h3A6]=8'h24; rom['h3A7]=8'h06;
    rom['h3A8]=8'h5B; rom['h3A9]=8'h5D; rom['h3AA]=8'h47; rom['h3AB]=8'hFD;
    rom['h3AC]=8'h20; rom['h3AD]=8'h04; rom['h3AE]=8'h48; rom['h3AF]=8'h6B;
    rom['h3B0]=8'h22; rom['h3B1]=8'h04; rom['h3B2]=8'h44; rom['h3B3]=8'h30;
    rom['h3B4]=8'h22; rom['h3B5]=8'h04; rom['h3B6]=8'h44; rom['h3B7]=8'h36;
    rom['h3B8]=8'h24; rom['h3B9]=8'h04; rom['h3BA]=8'h44; rom['h3BB]=8'h3C;
    rom['h3BC]=8'h20; rom['h3BD]=8'h00; rom['h3BE]=8'h58; rom['h3BF]=8'h11;
    rom['h3C0]=8'hA3; rom['h3C1]=8'hF4; rom['h3C2]=8'hB3; rom['h3C3]=8'hA2;
    rom['h3C4]=8'hF4; rom['h3C5]=8'hB2; rom['h3C6]=8'h47; rom['h3C7]=8'hF1;
    rom['h3C8]=8'hC0; rom['h3C9]=8'h5B; rom['h3CA]=8'h5D; rom['h3CB]=8'h24;
    rom['h3CC]=8'h18; rom['h3CD]=8'h57; rom['h3CE]=8'hFD; rom['h3CF]=8'h5B;
    rom['h3D0]=8'h5D; rom['h3D1]=8'h24; rom['h3D2]=8'h1A; rom['h3D3]=8'h47;
    rom['h3D4]=8'hFD; rom['h3D5]=8'h5B; rom['h3D6]=8'h5D; rom['h3D7]=8'h24;
    rom['h3D8]=8'h1C; rom['h3D9]=8'h57; rom['h3DA]=8'hFD; rom['h3DB]=8'h5B;
    rom['h3DC]=8'h5D; rom['h3DD]=8'h24; rom['h3DE]=8'h1E; rom['h3DF]=8'h57;
    rom['h3E0]=8'hFD; rom['h3E1]=8'h2E; rom['h3E2]=8'h00; rom['h3E3]=8'h58;
    rom['h3E4]=8'h09; rom['h3E5]=8'h20; rom['h3E6]=8'h1C; rom['h3E7]=8'h4B;
    rom['h3E8]=8'h81; rom['h3E9]=8'h20; rom['h3EA]=8'h18; rom['h3EB]=8'h48;
    rom['h3EC]=8'h5B; rom['h3ED]=8'h20; rom['h3EE]=8'h04; rom['h3EF]=8'h5B;
    rom['h3F0]=8'h5D; rom['h3F1]=8'h58; rom['h3F2]=8'h6B; rom['h3F3]=8'h5C;
    rom['h3F4]=8'hBF; rom['h3F5]=8'h5B; rom['h3F6]=8'h81; rom['h3F7]=8'h46;
    rom['h3F8]=8'hA6; rom['h3F9]=8'h20; rom['h3FA]=8'h04; rom['h3FB]=8'h5B;
    rom['h3FC]=8'h5D; rom['h3FD]=8'h58; rom['h3FE]=8'h6B; rom['h3FF]=8'h5C;
    rom['h400]=8'hCA; rom['h401]=8'h5B; rom['h402]=8'h81; rom['h403]=8'h46;
    rom['h404]=8'hA6; rom['h405]=8'h5B; rom['h406]=8'h5D; rom['h407]=8'h20;
    rom['h408]=8'h04; rom['h409]=8'h4B; rom['h40A]=8'h81; rom['h40B]=8'h46;
    rom['h40C]=8'h97; rom['h40D]=8'hC0; rom['h40E]=8'h20; rom['h40F]=8'h04;
    rom['h410]=8'h22; rom['h411]=8'h18; rom['h412]=8'h58; rom['h413]=8'hA0;
    rom['h414]=8'h46; rom['h415]=8'h8C; rom['h416]=8'h5B; rom['h417]=8'h5D;
    rom['h418]=8'h24; rom['h419]=8'h1C; rom['h41A]=8'h57; rom['h41B]=8'hFD;
    rom['h41C]=8'h5B; rom['h41D]=8'h5D; rom['h41E]=8'h24; rom['h41F]=8'h1E;
    rom['h420]=8'h57; rom['h421]=8'hFD; rom['h422]=8'h20; rom['h423]=8'h1C;
    rom['h424]=8'h5B; rom['h425]=8'h5D; rom['h426]=8'h24; rom['h427]=8'h00;
    rom['h428]=8'h47; rom['h429]=8'hFD; rom['h42A]=8'h20; rom['h42B]=8'h18;
    rom['h42C]=8'h48; rom['h42D]=8'h6B; rom['h42E]=8'h22; rom['h42F]=8'h00;
    rom['h430]=8'h57; rom['h431]=8'hAD; rom['h432]=8'h46; rom['h433]=8'hA4;
    rom['h434]=8'h22; rom['h435]=8'h00; rom['h436]=8'h57; rom['h437]=8'hBD;
    rom['h438]=8'h46; rom['h439]=8'hA4; rom['h43A]=8'h24; rom['h43B]=8'h00;
    rom['h43C]=8'h5B; rom['h43D]=8'h5D; rom['h43E]=8'h47; rom['h43F]=8'hFD;
    rom['h440]=8'h56; rom['h441]=8'h40; rom['h442]=8'hF3; rom['h443]=8'h46;
    rom['h444]=8'h8C; rom['h445]=8'h56; rom['h446]=8'h2D; rom['h447]=8'h44;
    rom['h448]=8'h8C; rom['h449]=8'h24; rom['h44A]=8'h0E; rom['h44B]=8'h26;
    rom['h44C]=8'h0C; rom['h44D]=8'h45; rom['h44E]=8'hC6; rom['h44F]=8'h56;
    rom['h450]=8'h2D; rom['h451]=8'h14; rom['h452]=8'h5F; rom['h453]=8'h58;
    rom['h454]=8'h5B; rom['h455]=8'h58; rom['h456]=8'h5B; rom['h457]=8'hC0;
    rom['h458]=8'h1C; rom['h459]=8'h5F; rom['h45A]=8'h58; rom['h45B]=8'h5B;
    rom['h45C]=8'h58; rom['h45D]=8'h5B; rom['h45E]=8'hC0; rom['h45F]=8'h5B;
    rom['h460]=8'h5D; rom['h461]=8'hA2; rom['h462]=8'hB6; rom['h463]=8'hA3;
    rom['h464]=8'hB7; rom['h465]=8'h5B; rom['h466]=8'h5D; rom['h467]=8'hA2;
    rom['h468]=8'hB4; rom['h469]=8'hA3; rom['h46A]=8'hB5; rom['h46B]=8'h47;
    rom['h46C]=8'h96; rom['h46D]=8'h56; rom['h46E]=8'h2D; rom['h46F]=8'h44;
    rom['h470]=8'hA3; rom['h471]=8'h24; rom['h472]=8'h0E; rom['h473]=8'h26;
    rom['h474]=8'h0C; rom['h475]=8'h45; rom['h476]=8'hDD; rom['h477]=8'h5B;
    rom['h478]=8'h5D; rom['h479]=8'h20; rom['h47A]=8'h00; rom['h47B]=8'h57;
    rom['h47C]=8'h9C; rom['h47D]=8'h56; rom['h47E]=8'h8C; rom['h47F]=8'h46;
    rom['h480]=8'hA0; rom['h481]=8'h24; rom['h482]=8'h00; rom['h483]=8'h26;
    rom['h484]=8'h00; rom['h485]=8'h44; rom['h486]=8'hB6; rom['h487]=8'h56;
    rom['h488]=8'h2D; rom['h489]=8'h1C; rom['h48A]=8'h8F; rom['h48B]=8'hC0;
    rom['h48C]=8'h14; rom['h48D]=8'h8F; rom['h48E]=8'hC0; rom['h48F]=8'h24;
    rom['h490]=8'h16; rom['h491]=8'h26; rom['h492]=8'h14; rom['h493]=8'h45;
    rom['h494]=8'hC6; rom['h495]=8'h56; rom['h496]=8'h2D; rom['h497]=8'h44;
    rom['h498]=8'h58; rom['h499]=8'hC0; rom['h49A]=8'h56; rom['h49B]=8'h2D;
    rom['h49C]=8'h1C; rom['h49D]=8'hAA; rom['h49E]=8'h58; rom['h49F]=8'h5B;
    rom['h4A0]=8'h58; rom['h4A1]=8'h5B; rom['h4A2]=8'hC0; rom['h4A3]=8'h14;
    rom['h4A4]=8'hAA; rom['h4A5]=8'h58; rom['h4A6]=8'h5B; rom['h4A7]=8'h58;
    rom['h4A8]=8'h5B; rom['h4A9]=8'hC0; rom['h4AA]=8'h5B; rom['h4AB]=8'h5D;
    rom['h4AC]=8'hA2; rom['h4AD]=8'hB6; rom['h4AE]=8'hA3; rom['h4AF]=8'hB7;
    rom['h4B0]=8'h5B; rom['h4B1]=8'h5D; rom['h4B2]=8'hA2; rom['h4B3]=8'hB4;
    rom['h4B4]=8'hA3; rom['h4B5]=8'hB5; rom['h4B6]=8'h22; rom['h4B7]=8'h1C;
    rom['h4B8]=8'h57; rom['h4B9]=8'h76; rom['h4BA]=8'h57; rom['h4BB]=8'h96;
    rom['h4BC]=8'h24; rom['h4BD]=8'h1E; rom['h4BE]=8'h26; rom['h4BF]=8'h1C;
    rom['h4C0]=8'h45; rom['h4C1]=8'hDD; rom['h4C2]=8'h5B; rom['h4C3]=8'h5D;
    rom['h4C4]=8'h20; rom['h4C5]=8'h00; rom['h4C6]=8'h56; rom['h4C7]=8'h40;
    rom['h4C8]=8'h1A; rom['h4C9]=8'hD3; rom['h4CA]=8'h5C; rom['h4CB]=8'hBF;
    rom['h4CC]=8'h1A; rom['h4CD]=8'hD3; rom['h4CE]=8'h57; rom['h4CF]=8'h9C;
    rom['h4D0]=8'hFA; rom['h4D1]=8'h44; rom['h4D2]=8'hD5; rom['h4D3]=8'h57;
    rom['h4D4]=8'h9C; rom['h4D5]=8'h56; rom['h4D6]=8'h8C; rom['h4D7]=8'h46;
    rom['h4D8]=8'hA0; rom['h4D9]=8'h24; rom['h4DA]=8'h00; rom['h4DB]=8'h26;
    rom['h4DC]=8'h08; rom['h4DD]=8'h44; rom['h4DE]=8'hB6; rom['h4DF]=8'h56;
    rom['h4E0]=8'h40; rom['h4E1]=8'h44; rom['h4E2]=8'h8C; rom['h4E3]=8'h24;
    rom['h4E4]=8'h0A; rom['h4E5]=8'h26; rom['h4E6]=8'h08; rom['h4E7]=8'h45;
    rom['h4E8]=8'hC6; rom['h4E9]=8'h56; rom['h4EA]=8'h40; rom['h4EB]=8'h44;
    rom['h4EC]=8'h51; rom['h4ED]=8'h5B; rom['h4EE]=8'h5D; rom['h4EF]=8'h49;
    rom['h4F0]=8'h69; rom['h4F1]=8'h56; rom['h4F2]=8'h40; rom['h4F3]=8'h44;
    rom['h4F4]=8'hA3; rom['h4F5]=8'h24; rom['h4F6]=8'h0A; rom['h4F7]=8'h26;
    rom['h4F8]=8'h08; rom['h4F9]=8'h45; rom['h4FA]=8'hDD; rom['h4FB]=8'h5B;
    rom['h4FC]=8'h5D; rom['h4FD]=8'h20; rom['h4FE]=8'h00; rom['h4FF]=8'h57;
    rom['h500]=8'hCD; rom['h501]=8'h56; rom['h502]=8'h8C; rom['h503]=8'h46;
    rom['h504]=8'hA0; rom['h505]=8'h24; rom['h506]=8'h00; rom['h507]=8'h26;
    rom['h508]=8'h10; rom['h509]=8'h44; rom['h50A]=8'hB6; rom['h50B]=8'h56;
    rom['h50C]=8'h40; rom['h50D]=8'h44; rom['h50E]=8'h89; rom['h50F]=8'hC0;
    rom['h510]=8'h56; rom['h511]=8'h40; rom['h512]=8'h44; rom['h513]=8'h58;
    rom['h514]=8'h5B; rom['h515]=8'h5D; rom['h516]=8'h49; rom['h517]=8'h81;
    rom['h518]=8'h56; rom['h519]=8'h40; rom['h51A]=8'h44; rom['h51B]=8'h9C;
    rom['h51C]=8'hC0; rom['h51D]=8'h5B; rom['h51E]=8'h5D; rom['h51F]=8'h56;
    rom['h520]=8'h40; rom['h521]=8'h14; rom['h522]=8'h25; rom['h523]=8'h5C;
    rom['h524]=8'hBF; rom['h525]=8'h20; rom['h526]=8'h00; rom['h527]=8'h57;
    rom['h528]=8'hCD; rom['h529]=8'h56; rom['h52A]=8'h8C; rom['h52B]=8'h46;
    rom['h52C]=8'hA0; rom['h52D]=8'h24; rom['h52E]=8'h00; rom['h52F]=8'h26;
    rom['h530]=8'h18; rom['h531]=8'h44; rom['h532]=8'hB6; rom['h533]=8'h56;
    rom['h534]=8'h7C; rom['h535]=8'h44; rom['h536]=8'h8C; rom['h537]=8'h24;
    rom['h538]=8'h06; rom['h539]=8'h26; rom['h53A]=8'h04; rom['h53B]=8'h45;
    rom['h53C]=8'hC6; rom['h53D]=8'h56; rom['h53E]=8'h7C; rom['h53F]=8'h44;
    rom['h540]=8'h51; rom['h541]=8'h24; rom['h542]=8'h1E; rom['h543]=8'h26;
    rom['h544]=8'h1C; rom['h545]=8'h20; rom['h546]=8'h18; rom['h547]=8'h5B;
    rom['h548]=8'h5D; rom['h549]=8'h57; rom['h54A]=8'hF7; rom['h54B]=8'h5B;
    rom['h54C]=8'h5D; rom['h54D]=8'h57; rom['h54E]=8'hFD; rom['h54F]=8'h24;
    rom['h550]=8'h06; rom['h551]=8'h26; rom['h552]=8'h04; rom['h553]=8'h58;
    rom['h554]=8'h1D; rom['h555]=8'h58; rom['h556]=8'h6B; rom['h557]=8'h5B;
    rom['h558]=8'h81; rom['h559]=8'h58; rom['h55A]=8'h23; rom['h55B]=8'h58;
    rom['h55C]=8'h6B; rom['h55D]=8'h5B; rom['h55E]=8'h81; rom['h55F]=8'h2C;
    rom['h560]=8'h04; rom['h561]=8'h2E; rom['h562]=8'h1C; rom['h563]=8'h48;
    rom['h564]=8'h50; rom['h565]=8'h56; rom['h566]=8'h7C; rom['h567]=8'h44;
    rom['h568]=8'hA3; rom['h569]=8'h24; rom['h56A]=8'h06; rom['h56B]=8'h26;
    rom['h56C]=8'h04; rom['h56D]=8'h45; rom['h56E]=8'hDD; rom['h56F]=8'h5B;
    rom['h570]=8'h5D; rom['h571]=8'hA2; rom['h572]=8'hB4; rom['h573]=8'hA3;
    rom['h574]=8'hB5; rom['h575]=8'h20; rom['h576]=8'h00; rom['h577]=8'h58;
    rom['h578]=8'h11; rom['h579]=8'h56; rom['h57A]=8'hB5; rom['h57B]=8'h57;
    rom['h57C]=8'hF1; rom['h57D]=8'h56; rom['h57E]=8'h8E; rom['h57F]=8'h46;
    rom['h580]=8'hA0; rom['h581]=8'h24; rom['h582]=8'h00; rom['h583]=8'h26;
    rom['h584]=8'h20; rom['h585]=8'h44; rom['h586]=8'hB6; rom['h587]=8'h56;
    rom['h588]=8'h7C; rom['h589]=8'h44; rom['h58A]=8'h89; rom['h58B]=8'h22;
    rom['h58C]=8'h04; rom['h58D]=8'h47; rom['h58E]=8'h6C; rom['h58F]=8'h56;
    rom['h590]=8'h7C; rom['h591]=8'h44; rom['h592]=8'h58; rom['h593]=8'h20;
    rom['h594]=8'h1C; rom['h595]=8'h22; rom['h596]=8'h04; rom['h597]=8'h57;
    rom['h598]=8'h6C; rom['h599]=8'h20; rom['h59A]=8'h08; rom['h59B]=8'h57;
    rom['h59C]=8'h76; rom['h59D]=8'h22; rom['h59E]=8'h1C; rom['h59F]=8'h47;
    rom['h5A0]=8'h6C; rom['h5A1]=8'h56; rom['h5A2]=8'h7C; rom['h5A3]=8'h44;
    rom['h5A4]=8'h9C; rom['h5A5]=8'hC0; rom['h5A6]=8'h5B; rom['h5A7]=8'h5D;
    rom['h5A8]=8'hA2; rom['h5A9]=8'hB4; rom['h5AA]=8'hA3; rom['h5AB]=8'hB5;
    rom['h5AC]=8'h20; rom['h5AD]=8'h00; rom['h5AE]=8'h58; rom['h5AF]=8'h11;
    rom['h5B0]=8'h56; rom['h5B1]=8'hC6; rom['h5B2]=8'h57; rom['h5B3]=8'hF1;
    rom['h5B4]=8'h56; rom['h5B5]=8'h8E; rom['h5B6]=8'h46; rom['h5B7]=8'hA0;
    rom['h5B8]=8'h24; rom['h5B9]=8'h00; rom['h5BA]=8'h26; rom['h5BB]=8'h28;
    rom['h5BC]=8'h44; rom['h5BD]=8'hB6; rom['h5BE]=8'h56; rom['h5BF]=8'h37;
    rom['h5C0]=8'h44; rom['h5C1]=8'h8C; rom['h5C2]=8'h24; rom['h5C3]=8'h00;
    rom['h5C4]=8'h26; rom['h5C5]=8'h10; rom['h5C6]=8'h20; rom['h5C7]=8'h18;
    rom['h5C8]=8'h5B; rom['h5C9]=8'h5D; rom['h5CA]=8'h57; rom['h5CB]=8'hF7;
    rom['h5CC]=8'h5B; rom['h5CD]=8'h5D; rom['h5CE]=8'h47; rom['h5CF]=8'hFD;
    rom['h5D0]=8'h56; rom['h5D1]=8'h37; rom['h5D2]=8'h44; rom['h5D3]=8'h51;
    rom['h5D4]=8'hC0; rom['h5D5]=8'h56; rom['h5D6]=8'h37; rom['h5D7]=8'h44;
    rom['h5D8]=8'hA3; rom['h5D9]=8'h24; rom['h5DA]=8'h00; rom['h5DB]=8'h26;
    rom['h5DC]=8'h10; rom['h5DD]=8'h20; rom['h5DE]=8'h18; rom['h5DF]=8'h58;
    rom['h5E0]=8'h1D; rom['h5E1]=8'h58; rom['h5E2]=8'h6B; rom['h5E3]=8'h5B;
    rom['h5E4]=8'h81; rom['h5E5]=8'h58; rom['h5E6]=8'h23; rom['h5E7]=8'h58;
    rom['h5E8]=8'h6B; rom['h5E9]=8'h4B; rom['h5EA]=8'h81; rom['h5EB]=8'h5B;
    rom['h5EC]=8'h5D; rom['h5ED]=8'hA2; rom['h5EE]=8'hB4; rom['h5EF]=8'hA3;
    rom['h5F0]=8'hB5; rom['h5F1]=8'h20; rom['h5F2]=8'h00; rom['h5F3]=8'h58;
    rom['h5F4]=8'h11; rom['h5F5]=8'h56; rom['h5F6]=8'hD7; rom['h5F7]=8'h57;
    rom['h5F8]=8'hF1; rom['h5F9]=8'h56; rom['h5FA]=8'h8E; rom['h5FB]=8'h46;
    rom['h5FC]=8'hA0; rom['h5FD]=8'h24; rom['h5FE]=8'h00; rom['h5FF]=8'h26;
    rom['h600]=8'h30; rom['h601]=8'h44; rom['h602]=8'hB6; rom['h603]=8'h56;
    rom['h604]=8'h37; rom['h605]=8'h44; rom['h606]=8'h89; rom['h607]=8'h2C;
    rom['h608]=8'h18; rom['h609]=8'h2E; rom['h60A]=8'h04; rom['h60B]=8'h48;
    rom['h60C]=8'h50; rom['h60D]=8'h56; rom['h60E]=8'h37; rom['h60F]=8'h44;
    rom['h610]=8'h58; rom['h611]=8'hC0; rom['h612]=8'h56; rom['h613]=8'h37;
    rom['h614]=8'h44; rom['h615]=8'h9C; rom['h616]=8'hC0; rom['h617]=8'h5B;
    rom['h618]=8'h5D; rom['h619]=8'h2C; rom['h61A]=8'h12; rom['h61B]=8'h2E;
    rom['h61C]=8'h00; rom['h61D]=8'h57; rom['h61E]=8'hE6; rom['h61F]=8'h20;
    rom['h620]=8'h12; rom['h621]=8'h57; rom['h622]=8'hCD; rom['h623]=8'h56;
    rom['h624]=8'h8C; rom['h625]=8'h46; rom['h626]=8'hA0; rom['h627]=8'h24;
    rom['h628]=8'h00; rom['h629]=8'h26; rom['h62A]=8'h38; rom['h62B]=8'h44;
    rom['h62C]=8'hB6; rom['h62D]=8'h2E; rom['h62E]=8'h11; rom['h62F]=8'h2F;
    rom['h630]=8'hE9; rom['h631]=8'hF5; rom['h632]=8'hF5; rom['h633]=8'h12;
    rom['h634]=8'h36; rom['h635]=8'hC0; rom['h636]=8'hC1; rom['h637]=8'h2E;
    rom['h638]=8'h11; rom['h639]=8'h2F; rom['h63A]=8'hE9; rom['h63B]=8'hF5;
    rom['h63C]=8'h12; rom['h63D]=8'h3F; rom['h63E]=8'hC0; rom['h63F]=8'hC1;
    rom['h640]=8'h2E; rom['h641]=8'h10; rom['h642]=8'h2F; rom['h643]=8'hE9;
    rom['h644]=8'hF6; rom['h645]=8'h12; rom['h646]=8'h48; rom['h647]=8'hC0;
    rom['h648]=8'hC1; rom['h649]=8'hF0; rom['h64A]=8'hBA; rom['h64B]=8'hA2;
    rom['h64C]=8'hF5; rom['h64D]=8'h1A; rom['h64E]=8'h50; rom['h64F]=8'h6A;
    rom['h650]=8'hF5; rom['h651]=8'h1A; rom['h652]=8'h54; rom['h653]=8'h6A;
    rom['h654]=8'hF5; rom['h655]=8'h1A; rom['h656]=8'h58; rom['h657]=8'h6A;
    rom['h658]=8'hF5; rom['h659]=8'h1A; rom['h65A]=8'h5C; rom['h65B]=8'h6A;
    rom['h65C]=8'hA3; rom['h65D]=8'hF5; rom['h65E]=8'h1A; rom['h65F]=8'h61;
    rom['h660]=8'h6A; rom['h661]=8'hF5; rom['h662]=8'h1A; rom['h663]=8'h65;
    rom['h664]=8'h6A; rom['h665]=8'hF5; rom['h666]=8'h1A; rom['h667]=8'h69;
    rom['h668]=8'h6A; rom['h669]=8'hF5; rom['h66A]=8'h1A; rom['h66B]=8'h6D;
    rom['h66C]=8'h6A; rom['h66D]=8'h2E; rom['h66E]=8'h10; rom['h66F]=8'h2F;
    rom['h670]=8'hE9; rom['h671]=8'hF5; rom['h672]=8'hF5; rom['h673]=8'hE0;
    rom['h674]=8'hAA; rom['h675]=8'hF6; rom['h676]=8'hF3; rom['h677]=8'hE9;
    rom['h678]=8'hF6; rom['h679]=8'hF6; rom['h67A]=8'hE0; rom['h67B]=8'hC0;
    rom['h67C]=8'h22; rom['h67D]=8'h00; rom['h67E]=8'h58; rom['h67F]=8'h17;
    rom['h680]=8'h56; rom['h681]=8'h49; rom['h682]=8'h2E; rom['h683]=8'h10;
    rom['h684]=8'h2F; rom['h685]=8'hE9; rom['h686]=8'hF5; rom['h687]=8'hF5;
    rom['h688]=8'h1A; rom['h689]=8'h8B; rom['h68A]=8'hC1; rom['h68B]=8'hC0;
    rom['h68C]=8'h12; rom['h68D]=8'h97; rom['h68E]=8'h2E; rom['h68F]=8'h10;
    rom['h690]=8'h2F; rom['h691]=8'hE9; rom['h692]=8'hF6; rom['h693]=8'hF1;
    rom['h694]=8'hF5; rom['h695]=8'hE0; rom['h696]=8'hC0; rom['h697]=8'h2E;
    rom['h698]=8'h10; rom['h699]=8'h2F; rom['h69A]=8'hE9; rom['h69B]=8'hF6;
    rom['h69C]=8'hFA; rom['h69D]=8'hF5; rom['h69E]=8'hE0; rom['h69F]=8'hC0;
    rom['h6A0]=8'h58; rom['h6A1]=8'h11; rom['h6A2]=8'h46; rom['h6A3]=8'hA6;
    rom['h6A4]=8'h58; rom['h6A5]=8'h17; rom['h6A6]=8'hA2; rom['h6A7]=8'hF5;
    rom['h6A8]=8'hF7; rom['h6A9]=8'hBA; rom['h6AA]=8'h5D; rom['h6AB]=8'h34;
    rom['h6AC]=8'hF6; rom['h6AD]=8'hF3; rom['h6AE]=8'hAA; rom['h6AF]=8'hF6;
    rom['h6B0]=8'hF6; rom['h6B1]=8'h2E; rom['h6B2]=8'h11; rom['h6B3]=8'h2F;
    rom['h6B4]=8'hE0; rom['h6B5]=8'hA3; rom['h6B6]=8'hB6; rom['h6B7]=8'hA5;
    rom['h6B8]=8'hB7; rom['h6B9]=8'h56; rom['h6BA]=8'hE8; rom['h6BB]=8'hA6;
    rom['h6BC]=8'hB3; rom['h6BD]=8'hA2; rom['h6BE]=8'hB6; rom['h6BF]=8'hA4;
    rom['h6C0]=8'hB7; rom['h6C1]=8'h56; rom['h6C2]=8'hE8; rom['h6C3]=8'hA6;
    rom['h6C4]=8'hB2; rom['h6C5]=8'hC0; rom['h6C6]=8'hA3; rom['h6C7]=8'hB6;
    rom['h6C8]=8'hA5; rom['h6C9]=8'hB7; rom['h6CA]=8'h57; rom['h6CB]=8'h14;
    rom['h6CC]=8'hA6; rom['h6CD]=8'hB3; rom['h6CE]=8'hA2; rom['h6CF]=8'hB6;
    rom['h6D0]=8'hA4; rom['h6D1]=8'hB7; rom['h6D2]=8'h57; rom['h6D3]=8'h14;
    rom['h6D4]=8'hA6; rom['h6D5]=8'hB2; rom['h6D6]=8'hC0; rom['h6D7]=8'hA3;
    rom['h6D8]=8'hB6; rom['h6D9]=8'hA5; rom['h6DA]=8'hB7; rom['h6DB]=8'h57;
    rom['h6DC]=8'h40; rom['h6DD]=8'hA6; rom['h6DE]=8'hB3; rom['h6DF]=8'hA2;
    rom['h6E0]=8'hB6; rom['h6E1]=8'hA4; rom['h6E2]=8'hB7; rom['h6E3]=8'h57;
    rom['h6E4]=8'h40; rom['h6E5]=8'hA6; rom['h6E6]=8'hB2; rom['h6E7]=8'hC0;
    rom['h6E8]=8'hF0; rom['h6E9]=8'hA7; rom['h6EA]=8'hF6; rom['h6EB]=8'h12;
    rom['h6EC]=8'hF2; rom['h6ED]=8'hA6; rom['h6EE]=8'hF6; rom['h6EF]=8'hF1;
    rom['h6F0]=8'hF5; rom['h6F1]=8'hB6; rom['h6F2]=8'hA7; rom['h6F3]=8'hF6;
    rom['h6F4]=8'hF6; rom['h6F5]=8'h12; rom['h6F6]=8'hFE; rom['h6F7]=8'hA6;
    rom['h6F8]=8'hF6; rom['h6F9]=8'hF6; rom['h6FA]=8'hF1; rom['h6FB]=8'hF5;
    rom['h6FC]=8'hF5; rom['h6FD]=8'hB6; rom['h6FE]=8'hA7; rom['h6FF]=8'hF5;
    rom['h700]=8'hF5; rom['h701]=8'h12; rom['h702]=8'h0A; rom['h703]=8'hA6;
    rom['h704]=8'hF5; rom['h705]=8'hF5; rom['h706]=8'hF1; rom['h707]=8'hF6;
    rom['h708]=8'hF6; rom['h709]=8'hB6; rom['h70A]=8'hA7; rom['h70B]=8'hF5;
    rom['h70C]=8'h12; rom['h70D]=8'h13; rom['h70E]=8'hA6; rom['h70F]=8'hF5;
    rom['h710]=8'hF1; rom['h711]=8'hF6; rom['h712]=8'hB6; rom['h713]=8'hC0;
    rom['h714]=8'hF0; rom['h715]=8'hA7; rom['h716]=8'hF6; rom['h717]=8'h1A;
    rom['h718]=8'h1E; rom['h719]=8'hA6; rom['h71A]=8'hF6; rom['h71B]=8'hF3;
    rom['h71C]=8'hF5; rom['h71D]=8'hB6; rom['h71E]=8'hA7; rom['h71F]=8'hF6;
    rom['h720]=8'hF6; rom['h721]=8'h1A; rom['h722]=8'h2A; rom['h723]=8'hA6;
    rom['h724]=8'hF6; rom['h725]=8'hF6; rom['h726]=8'hF3; rom['h727]=8'hF5;
    rom['h728]=8'hF5; rom['h729]=8'hB6; rom['h72A]=8'hA7; rom['h72B]=8'hF5;
    rom['h72C]=8'hF5; rom['h72D]=8'h1A; rom['h72E]=8'h36; rom['h72F]=8'hA6;
    rom['h730]=8'hF5; rom['h731]=8'hF5; rom['h732]=8'hF3; rom['h733]=8'hF6;
    rom['h734]=8'hF6; rom['h735]=8'hB6; rom['h736]=8'hA7; rom['h737]=8'hF5;
    rom['h738]=8'h1A; rom['h739]=8'h3F; rom['h73A]=8'hA6; rom['h73B]=8'hF5;
    rom['h73C]=8'hF3; rom['h73D]=8'hF6; rom['h73E]=8'hB6; rom['h73F]=8'hC0;
    rom['h740]=8'hF0; rom['h741]=8'hA7; rom['h742]=8'hF6; rom['h743]=8'h1A;
    rom['h744]=8'h4A; rom['h745]=8'hA6; rom['h746]=8'hF6; rom['h747]=8'hFA;
    rom['h748]=8'hF5; rom['h749]=8'hB6; rom['h74A]=8'hA7; rom['h74B]=8'hF6;
    rom['h74C]=8'hF6; rom['h74D]=8'h1A; rom['h74E]=8'h56; rom['h74F]=8'hA6;
    rom['h750]=8'hF6; rom['h751]=8'hF6; rom['h752]=8'hFA; rom['h753]=8'hF5;
    rom['h754]=8'hF5; rom['h755]=8'hB6; rom['h756]=8'hA7; rom['h757]=8'hF5;
    rom['h758]=8'hF5; rom['h759]=8'h1A; rom['h75A]=8'h62; rom['h75B]=8'hA6;
    rom['h75C]=8'hF5; rom['h75D]=8'hF5; rom['h75E]=8'hFA; rom['h75F]=8'hF6;
    rom['h760]=8'hF6; rom['h761]=8'hB6; rom['h762]=8'hA7; rom['h763]=8'hF5;
    rom['h764]=8'h1A; rom['h765]=8'h6B; rom['h766]=8'hA6; rom['h767]=8'hF5;
    rom['h768]=8'hFA; rom['h769]=8'hF6; rom['h76A]=8'hB6; rom['h76B]=8'hC0;
    rom['h76C]=8'hA0; rom['h76D]=8'hBC; rom['h76E]=8'hA1; rom['h76F]=8'hBD;
    rom['h770]=8'hA2; rom['h771]=8'hBE; rom['h772]=8'hA3; rom['h773]=8'hBF;
    rom['h774]=8'h48; rom['h775]=8'h50; rom['h776]=8'hA2; rom['h777]=8'hBC;
    rom['h778]=8'hA3; rom['h779]=8'hBD; rom['h77A]=8'hA0; rom['h77B]=8'hBE;
    rom['h77C]=8'hA1; rom['h77D]=8'hBF; rom['h77E]=8'h48; rom['h77F]=8'h50;
    rom['h780]=8'h2F; rom['h781]=8'hA7; rom['h782]=8'hE0; rom['h783]=8'h6F;
    rom['h784]=8'h2F; rom['h785]=8'hA6; rom['h786]=8'hE0; rom['h787]=8'h6F;
    rom['h788]=8'h2F; rom['h789]=8'hA5; rom['h78A]=8'hE0; rom['h78B]=8'h6F;
    rom['h78C]=8'h2F; rom['h78D]=8'hA4; rom['h78E]=8'hE0; rom['h78F]=8'hC0;
    rom['h790]=8'hA2; rom['h791]=8'hBE; rom['h792]=8'hA3; rom['h793]=8'hBF;
    rom['h794]=8'h47; rom['h795]=8'h80; rom['h796]=8'hA0; rom['h797]=8'hBE;
    rom['h798]=8'hA1; rom['h799]=8'hBF; rom['h79A]=8'h47; rom['h79B]=8'h80;
    rom['h79C]=8'hA0; rom['h79D]=8'hBE; rom['h79E]=8'hA1; rom['h79F]=8'hBF;
    rom['h7A0]=8'h2F; rom['h7A1]=8'hE9; rom['h7A2]=8'hA3; rom['h7A3]=8'hF1;
    rom['h7A4]=8'hEB; rom['h7A5]=8'hE0; rom['h7A6]=8'h6F; rom['h7A7]=8'h2F;
    rom['h7A8]=8'hE9; rom['h7A9]=8'hA2; rom['h7AA]=8'hEB; rom['h7AB]=8'hE0;
    rom['h7AC]=8'hC0; rom['h7AD]=8'hA2; rom['h7AE]=8'hBE; rom['h7AF]=8'hA3;
    rom['h7B0]=8'hBF; rom['h7B1]=8'h2F; rom['h7B2]=8'hE9; rom['h7B3]=8'hF2;
    rom['h7B4]=8'hE0; rom['h7B5]=8'h1C; rom['h7B6]=8'hBC; rom['h7B7]=8'h6F;
    rom['h7B8]=8'h2F; rom['h7B9]=8'hE9; rom['h7BA]=8'hF2; rom['h7BB]=8'hE0;
    rom['h7BC]=8'hC0; rom['h7BD]=8'hA2; rom['h7BE]=8'hBE; rom['h7BF]=8'hA3;
    rom['h7C0]=8'hBF; rom['h7C1]=8'h2F; rom['h7C2]=8'hE9; rom['h7C3]=8'hF8;
    rom['h7C4]=8'hE0; rom['h7C5]=8'h12; rom['h7C6]=8'hCC; rom['h7C7]=8'h6F;
    rom['h7C8]=8'h2F; rom['h7C9]=8'hE9; rom['h7CA]=8'hF8; rom['h7CB]=8'hE0;
    rom['h7CC]=8'hC0; rom['h7CD]=8'hA0; rom['h7CE]=8'hBE; rom['h7CF]=8'hA1;
    rom['h7D0]=8'hBF; rom['h7D1]=8'h2F; rom['h7D2]=8'hE9; rom['h7D3]=8'hF1;
    rom['h7D4]=8'h93; rom['h7D5]=8'hE0; rom['h7D6]=8'hF3; rom['h7D7]=8'h6F;
    rom['h7D8]=8'h2F; rom['h7D9]=8'hE9; rom['h7DA]=8'h92; rom['h7DB]=8'hE0;
    rom['h7DC]=8'hF3; rom['h7DD]=8'hC0; rom['h7DE]=8'hA0; rom['h7DF]=8'hBC;
    rom['h7E0]=8'hA1; rom['h7E1]=8'hBD; rom['h7E2]=8'hA2; rom['h7E3]=8'hBE;
    rom['h7E4]=8'hA3; rom['h7E5]=8'hBF; rom['h7E6]=8'h2F; rom['h7E7]=8'hE9;
    rom['h7E8]=8'h2D; rom['h7E9]=8'hE0; rom['h7EA]=8'h6F; rom['h7EB]=8'h6D;
    rom['h7EC]=8'h2F; rom['h7ED]=8'hE9; rom['h7EE]=8'h2D; rom['h7EF]=8'hE0;
    rom['h7F0]=8'hC0; rom['h7F1]=8'hA0; rom['h7F2]=8'hBE; rom['h7F3]=8'hA1;
    rom['h7F4]=8'hBF; rom['h7F5]=8'h48; rom['h7F6]=8'h01; rom['h7F7]=8'hA6;
    rom['h7F8]=8'hBE; rom['h7F9]=8'hA7; rom['h7FA]=8'hBF; rom['h7FB]=8'h48;
    rom['h7FC]=8'h01; rom['h7FD]=8'hA4; rom['h7FE]=8'hBE; rom['h7FF]=8'hA5;
    rom['h800]=8'hBF; rom['h801]=8'h2F; rom['h802]=8'hA3; rom['h803]=8'hE0;
    rom['h804]=8'h6F; rom['h805]=8'h2F; rom['h806]=8'hA2; rom['h807]=8'hE0;
    rom['h808]=8'hC0; rom['h809]=8'h2F; rom['h80A]=8'hE9; rom['h80B]=8'hB3;
    rom['h80C]=8'h6F; rom['h80D]=8'h2F; rom['h80E]=8'hE9; rom['h80F]=8'hB2;
    rom['h810]=8'hC0; rom['h811]=8'hA0; rom['h812]=8'hBE; rom['h813]=8'hA1;
    rom['h814]=8'hBF; rom['h815]=8'h48; rom['h816]=8'h09; rom['h817]=8'hA2;
    rom['h818]=8'hBE; rom['h819]=8'hA3; rom['h81A]=8'hBF; rom['h81B]=8'h48;
    rom['h81C]=8'h09; rom['h81D]=8'hA4; rom['h81E]=8'hBE; rom['h81F]=8'hA5;
    rom['h820]=8'hBF; rom['h821]=8'h48; rom['h822]=8'h09; rom['h823]=8'hA6;
    rom['h824]=8'hBE; rom['h825]=8'hA7; rom['h826]=8'hBF; rom['h827]=8'h48;
    rom['h828]=8'h09; rom['h829]=8'h5B; rom['h82A]=8'h00; rom['h82B]=8'hA6;
    rom['h82C]=8'hB0; rom['h82D]=8'hA7; rom['h82E]=8'hB1; rom['h82F]=8'h5B;
    rom['h830]=8'h00; rom['h831]=8'h5B; rom['h832]=8'h12; rom['h833]=8'h5B;
    rom['h834]=8'h24; rom['h835]=8'h58; rom['h836]=8'hB5; rom['h837]=8'hA4;
    rom['h838]=8'h5C; rom['h839]=8'hB4; rom['h83A]=8'hA5; rom['h83B]=8'h5C;
    rom['h83C]=8'hB4; rom['h83D]=8'hA6; rom['h83E]=8'h5C; rom['h83F]=8'hB4;
    rom['h840]=8'hA7; rom['h841]=8'h5C; rom['h842]=8'hB4; rom['h843]=8'h5B;
    rom['h844]=8'h50; rom['h845]=8'h5B; rom['h846]=8'h43; rom['h847]=8'h5B;
    rom['h848]=8'h36; rom['h849]=8'hA0; rom['h84A]=8'hB6; rom['h84B]=8'hA1;
    rom['h84C]=8'hB7; rom['h84D]=8'h5B; rom['h84E]=8'h36; rom['h84F]=8'hC0;
    rom['h850]=8'hDC; rom['h851]=8'hBB; rom['h852]=8'h2F; rom['h853]=8'hE9;
    rom['h854]=8'h2D; rom['h855]=8'hE0; rom['h856]=8'h6F; rom['h857]=8'h6D;
    rom['h858]=8'h7B; rom['h859]=8'h52; rom['h85A]=8'hC0; rom['h85B]=8'hA1;
    rom['h85C]=8'hBF; rom['h85D]=8'hDC; rom['h85E]=8'hBE; rom['h85F]=8'h21;
    rom['h860]=8'hE9; rom['h861]=8'hF2; rom['h862]=8'hE0; rom['h863]=8'h1C;
    rom['h864]=8'h68; rom['h865]=8'h61; rom['h866]=8'h7E; rom['h867]=8'h5F;
    rom['h868]=8'hAF; rom['h869]=8'hB1; rom['h86A]=8'hC0; rom['h86B]=8'hA1;
    rom['h86C]=8'hBF; rom['h86D]=8'hDC; rom['h86E]=8'hBE; rom['h86F]=8'hF1;
    rom['h870]=8'h21; rom['h871]=8'hE9; rom['h872]=8'hF8; rom['h873]=8'hE0;
    rom['h874]=8'h12; rom['h875]=8'h79; rom['h876]=8'h61; rom['h877]=8'h7E;
    rom['h878]=8'h70; rom['h879]=8'hAF; rom['h87A]=8'hB1; rom['h87B]=8'hC0;
    rom['h87C]=8'hA1; rom['h87D]=8'hBF; rom['h87E]=8'hA3; rom['h87F]=8'hBD;
    rom['h880]=8'hF0; rom['h881]=8'hBC; rom['h882]=8'hDC; rom['h883]=8'hBE;
    rom['h884]=8'hFA; rom['h885]=8'hF3; rom['h886]=8'h21; rom['h887]=8'hE9;
    rom['h888]=8'h23; rom['h889]=8'hE8; rom['h88A]=8'h61; rom['h88B]=8'h63;
    rom['h88C]=8'hBB; rom['h88D]=8'hAB; rom['h88E]=8'h14; rom['h88F]=8'h92;
    rom['h890]=8'hD1; rom['h891]=8'hBC; rom['h892]=8'h7E; rom['h893]=8'h85;
    rom['h894]=8'hAB; rom['h895]=8'hF5; rom['h896]=8'hF3; rom['h897]=8'hAF;
    rom['h898]=8'hB1; rom['h899]=8'hAD; rom['h89A]=8'hB3; rom['h89B]=8'hAC;
    rom['h89C]=8'h14; rom['h89D]=8'h9F; rom['h89E]=8'hC1; rom['h89F]=8'hC0;
    rom['h8A0]=8'hA1; rom['h8A1]=8'hBF; rom['h8A2]=8'hA3; rom['h8A3]=8'hBD;
    rom['h8A4]=8'hDC; rom['h8A5]=8'hBE; rom['h8A6]=8'hF1; rom['h8A7]=8'h23;
    rom['h8A8]=8'hE9; rom['h8A9]=8'h21; rom['h8AA]=8'hEB; rom['h8AB]=8'hE0;
    rom['h8AC]=8'h61; rom['h8AD]=8'h63; rom['h8AE]=8'h7E; rom['h8AF]=8'hA7;
    rom['h8B0]=8'hAF; rom['h8B1]=8'hB1; rom['h8B2]=8'hAD; rom['h8B3]=8'hB3;
    rom['h8B4]=8'hC0; rom['h8B5]=8'hA2; rom['h8B6]=8'hBE; rom['h8B7]=8'hA3;
    rom['h8B8]=8'hBF; rom['h8B9]=8'h2F; rom['h8BA]=8'hE9; rom['h8BB]=8'hB7;
    rom['h8BC]=8'h6F; rom['h8BD]=8'h2F; rom['h8BE]=8'hE9; rom['h8BF]=8'hB6;
    rom['h8C0]=8'h6F; rom['h8C1]=8'h2F; rom['h8C2]=8'hE9; rom['h8C3]=8'hB5;
    rom['h8C4]=8'h6F; rom['h8C5]=8'h2F; rom['h8C6]=8'hE9; rom['h8C7]=8'hB4;
    rom['h8C8]=8'hC0; rom['h8C9]=8'h5B; rom['h8CA]=8'h12; rom['h8CB]=8'h5B;
    rom['h8CC]=8'h5D; rom['h8CD]=8'h5C; rom['h8CE]=8'hF0; rom['h8CF]=8'h1C;
    rom['h8D0]=8'hD4; rom['h8D1]=8'h5B; rom['h8D2]=8'h43; rom['h8D3]=8'hC1;
    rom['h8D4]=8'h24; rom['h8D5]=8'h00; rom['h8D6]=8'h26; rom['h8D7]=8'h00;
    rom['h8D8]=8'h5D; rom['h8D9]=8'h1B; rom['h8DA]=8'h5E; rom['h8DB]=8'h16;
    rom['h8DC]=8'hA3; rom['h8DD]=8'hB7; rom['h8DE]=8'h5B; rom['h8DF]=8'h5D;
    rom['h8E0]=8'h5C; rom['h8E1]=8'hF0; rom['h8E2]=8'h14; rom['h8E3]=8'hE6;
    rom['h8E4]=8'h48; rom['h8E5]=8'hD8; rom['h8E6]=8'h5B; rom['h8E7]=8'h43;
    rom['h8E8]=8'h47; rom['h8E9]=8'h90; rom['h8EA]=8'h20; rom['h8EB]=8'h87;
    rom['h8EC]=8'h5E; rom['h8ED]=8'h00; rom['h8EE]=8'h22; rom['h8EF]=8'h00;
    rom['h8F0]=8'h58; rom['h8F1]=8'h17; rom['h8F2]=8'h5C; rom['h8F3]=8'h85;
    rom['h8F4]=8'h5C; rom['h8F5]=8'h98; rom['h8F6]=8'h56; rom['h8F7]=8'h37;
    rom['h8F8]=8'h5C; rom['h8F9]=8'hB4; rom['h8FA]=8'h56; rom['h8FB]=8'h2D;
    rom['h8FC]=8'h5C; rom['h8FD]=8'hB4; rom['h8FE]=8'h56; rom['h8FF]=8'h40;
    rom['h900]=8'h5C; rom['h901]=8'hB4; rom['h902]=8'h5C; rom['h903]=8'h98;
    rom['h904]=8'h22; rom['h905]=8'h0C; rom['h906]=8'h58; rom['h907]=8'h29;
    rom['h908]=8'h5C; rom['h909]=8'h98; rom['h90A]=8'h22; rom['h90B]=8'h08;
    rom['h90C]=8'h58; rom['h90D]=8'h29; rom['h90E]=8'h5C; rom['h90F]=8'h98;
    rom['h910]=8'h22; rom['h911]=8'h04; rom['h912]=8'h58; rom['h913]=8'h29;
    rom['h914]=8'h5C; rom['h915]=8'h98; rom['h916]=8'h22; rom['h917]=8'h18;
    rom['h918]=8'h58; rom['h919]=8'h29; rom['h91A]=8'h5C; rom['h91B]=8'h98;
    rom['h91C]=8'h22; rom['h91D]=8'h14; rom['h91E]=8'h58; rom['h91F]=8'h29;
    rom['h920]=8'h5C; rom['h921]=8'h98; rom['h922]=8'h20; rom['h923]=8'h1C;
    rom['h924]=8'h22; rom['h925]=8'h14; rom['h926]=8'h57; rom['h927]=8'h6C;
    rom['h928]=8'h5B; rom['h929]=8'h5D; rom['h92A]=8'h5C; rom['h92B]=8'h85;
    rom['h92C]=8'h5C; rom['h92D]=8'h98; rom['h92E]=8'h5B; rom['h92F]=8'h5D;
    rom['h930]=8'h5C; rom['h931]=8'h85; rom['h932]=8'h5C; rom['h933]=8'h98;
    rom['h934]=8'h5B; rom['h935]=8'h5D; rom['h936]=8'h5C; rom['h937]=8'h85;
    rom['h938]=8'h5C; rom['h939]=8'h98; rom['h93A]=8'h20; rom['h93B]=8'h0C;
    rom['h93C]=8'h5B; rom['h93D]=8'h5D; rom['h93E]=8'h58; rom['h93F]=8'h6B;
    rom['h940]=8'h5C; rom['h941]=8'h85; rom['h942]=8'h5C; rom['h943]=8'h98;
    rom['h944]=8'h20; rom['h945]=8'h08; rom['h946]=8'h5B; rom['h947]=8'h5D;
    rom['h948]=8'h58; rom['h949]=8'h6B; rom['h94A]=8'h5C; rom['h94B]=8'h85;
    rom['h94C]=8'h5C; rom['h94D]=8'h98; rom['h94E]=8'h20; rom['h94F]=8'h04;
    rom['h950]=8'h5B; rom['h951]=8'h5D; rom['h952]=8'h58; rom['h953]=8'h6B;
    rom['h954]=8'h5C; rom['h955]=8'h85; rom['h956]=8'h5C; rom['h957]=8'h98;
    rom['h958]=8'h20; rom['h959]=8'h18; rom['h95A]=8'h5B; rom['h95B]=8'h5D;
    rom['h95C]=8'h5C; rom['h95D]=8'h85; rom['h95E]=8'h5C; rom['h95F]=8'h98;
    rom['h960]=8'h5B; rom['h961]=8'h5D; rom['h962]=8'h5C; rom['h963]=8'h85;
    rom['h964]=8'h58; rom['h965]=8'h6B; rom['h966]=8'h58; rom['h967]=8'h6B;
    rom['h968]=8'hC0; rom['h969]=8'h2E; rom['h96A]=8'h00; rom['h96B]=8'h5D;
    rom['h96C]=8'h27; rom['h96D]=8'h1C; rom['h96E]=8'h71; rom['h96F]=8'h49;
    rom['h970]=8'h7A; rom['h971]=8'h2E; rom['h972]=8'h01; rom['h973]=8'h5D;
    rom['h974]=8'h27; rom['h975]=8'h1C; rom['h976]=8'h79; rom['h977]=8'h49;
    rom['h978]=8'h80; rom['h979]=8'hC0; rom['h97A]=8'h22; rom['h97B]=8'h00;
    rom['h97C]=8'h58; rom['h97D]=8'h17; rom['h97E]=8'h4C; rom['h97F]=8'h5F;
    rom['h980]=8'hC0; rom['h981]=8'h2E; rom['h982]=8'h00; rom['h983]=8'h5D;
    rom['h984]=8'h27; rom['h985]=8'h1C; rom['h986]=8'h89; rom['h987]=8'h49;
    rom['h988]=8'h92; rom['h989]=8'h2E; rom['h98A]=8'h01; rom['h98B]=8'h5D;
    rom['h98C]=8'h27; rom['h98D]=8'h1C; rom['h98E]=8'h91; rom['h98F]=8'h49;
    rom['h990]=8'hB2; rom['h991]=8'hC0; rom['h992]=8'h2E; rom['h993]=8'h20;
    rom['h994]=8'h58; rom['h995]=8'h09; rom['h996]=8'h5D; rom['h997]=8'h34;
    rom['h998]=8'h1C; rom['h999]=8'h9C; rom['h99A]=8'h5C; rom['h99B]=8'h37;
    rom['h99C]=8'h2E; rom['h99D]=8'h1B; rom['h99E]=8'h5D; rom['h99F]=8'h27;
    rom['h9A0]=8'h14; rom['h9A1]=8'hAC; rom['h9A2]=8'h20; rom['h9A3]=8'h00;
    rom['h9A4]=8'h57; rom['h9A5]=8'hF1; rom['h9A6]=8'h2E; rom['h9A7]=8'h20;
    rom['h9A8]=8'h22; rom['h9A9]=8'h00; rom['h9AA]=8'h48; rom['h9AB]=8'h01;
    rom['h9AC]=8'h5C; rom['h9AD]=8'hA0; rom['h9AE]=8'h58; rom['h9AF]=8'hEA;
    rom['h9B0]=8'h40; rom['h9B1]=8'h2D; rom['h9B2]=8'h19; rom['h9B3]=8'hBC;
    rom['h9B4]=8'h11; rom['h9B5]=8'hB4; rom['h9B6]=8'h20; rom['h9B7]=8'h20;
    rom['h9B8]=8'h22; rom['h9B9]=8'h03; rom['h9BA]=8'h47; rom['h9BB]=8'hF1;
    rom['h9BC]=8'h20; rom['h9BD]=8'h00; rom['h9BE]=8'h22; rom['h9BF]=8'hFF;
    rom['h9C0]=8'h47; rom['h9C1]=8'hF1; rom['h9C2]=8'hFF; rom['h9C3]=8'hFF;
    rom['h9C4]=8'hFF; rom['h9C5]=8'hFF; rom['h9C6]=8'hFF; rom['h9C7]=8'hFF;
    rom['h9C8]=8'hFF; rom['h9C9]=8'hFF; rom['h9CA]=8'hFF; rom['h9CB]=8'hFF;
    rom['h9CC]=8'hFF; rom['h9CD]=8'hFF; rom['h9CE]=8'hFF; rom['h9CF]=8'hFF;
    rom['h9D0]=8'hFF; rom['h9D1]=8'hFF; rom['h9D2]=8'hFF; rom['h9D3]=8'hFF;
    rom['h9D4]=8'hFF; rom['h9D5]=8'hFF; rom['h9D6]=8'hFF; rom['h9D7]=8'hFF;
    rom['h9D8]=8'hFF; rom['h9D9]=8'hFF; rom['h9DA]=8'hFF; rom['h9DB]=8'hFF;
    rom['h9DC]=8'hFF; rom['h9DD]=8'hFF; rom['h9DE]=8'hFF; rom['h9DF]=8'hFF;
    rom['h9E0]=8'hFF; rom['h9E1]=8'hFF; rom['h9E2]=8'hFF; rom['h9E3]=8'hFF;
    rom['h9E4]=8'hFF; rom['h9E5]=8'hFF; rom['h9E6]=8'hFF; rom['h9E7]=8'hFF;
    rom['h9E8]=8'hFF; rom['h9E9]=8'hFF; rom['h9EA]=8'hFF; rom['h9EB]=8'hFF;
    rom['h9EC]=8'hFF; rom['h9ED]=8'hFF; rom['h9EE]=8'hFF; rom['h9EF]=8'h35;
    rom['h9F0]=8'h44; rom['h9F1]=8'h79; rom['h9F2]=8'h44; rom['h9F3]=8'hC4;
    rom['h9F4]=8'h44; rom['h9F5]=8'hFD; rom['h9F6]=8'h45; rom['h9F7]=8'h1F;
    rom['h9F8]=8'h45; rom['h9F9]=8'h71; rom['h9FA]=8'h45; rom['h9FB]=8'hA8;
    rom['h9FC]=8'h45; rom['h9FD]=8'hED; rom['h9FE]=8'h46; rom['h9FF]=8'h19;
    rom['hA00]=8'h33; rom['hA01]=8'h00; rom['hA02]=8'h42; rom['hA03]=8'h72;
    rom['hA04]=8'h42; rom['hA05]=8'h7E; rom['hA06]=8'h42; rom['hA07]=8'h86;
    rom['hA08]=8'h42; rom['hA09]=8'h8A; rom['hA0A]=8'h42; rom['hA0B]=8'h8E;
    rom['hA0C]=8'h42; rom['hA0D]=8'h92; rom['hA0E]=8'h42; rom['hA0F]=8'h96;
    rom['hA10]=8'h42; rom['hA11]=8'hA6; rom['hA12]=8'h42; rom['hA13]=8'hA7;
    rom['hA14]=8'h42; rom['hA15]=8'hAF; rom['hA16]=8'h42; rom['hA17]=8'hB9;
    rom['hA18]=8'h42; rom['hA19]=8'hBD; rom['hA1A]=8'h42; rom['hA1B]=8'hC1;
    rom['hA1C]=8'h42; rom['hA1D]=8'hC5; rom['hA1E]=8'h42; rom['hA1F]=8'hC9;
    rom['hA20]=8'h42; rom['hA21]=8'hD9; rom['hA22]=8'h42; rom['hA23]=8'hDA;
    rom['hA24]=8'h42; rom['hA25]=8'hE6; rom['hA26]=8'h42; rom['hA27]=8'hEE;
    rom['hA28]=8'h42; rom['hA29]=8'hF2; rom['hA2A]=8'h42; rom['hA2B]=8'hF6;
    rom['hA2C]=8'h42; rom['hA2D]=8'hFA; rom['hA2E]=8'h42; rom['hA2F]=8'hFE;
    rom['hA30]=8'h43; rom['hA31]=8'h0E; rom['hA32]=8'h43; rom['hA33]=8'h0F;
    rom['hA34]=8'h43; rom['hA35]=8'h17; rom['hA36]=8'h43; rom['hA37]=8'h21;
    rom['hA38]=8'h43; rom['hA39]=8'h25; rom['hA3A]=8'h43; rom['hA3B]=8'h29;
    rom['hA3C]=8'h43; rom['hA3D]=8'h2D; rom['hA3E]=8'h43; rom['hA3F]=8'h31;
    rom['hA40]=8'h43; rom['hA41]=8'h41; rom['hA42]=8'h43; rom['hA43]=8'h42;
    rom['hA44]=8'h43; rom['hA45]=8'h4E; rom['hA46]=8'h43; rom['hA47]=8'h6C;
    rom['hA48]=8'h43; rom['hA49]=8'h70; rom['hA4A]=8'h43; rom['hA4B]=8'h74;
    rom['hA4C]=8'h43; rom['hA4D]=8'h78; rom['hA4E]=8'h43; rom['hA4F]=8'h7C;
    rom['hA50]=8'h43; rom['hA51]=8'h89; rom['hA52]=8'h43; rom['hA53]=8'h8A;
    rom['hA54]=8'h43; rom['hA55]=8'h92; rom['hA56]=8'h43; rom['hA57]=8'hAC;
    rom['hA58]=8'h43; rom['hA59]=8'hB0; rom['hA5A]=8'h43; rom['hA5B]=8'hB4;
    rom['hA5C]=8'h43; rom['hA5D]=8'hB8; rom['hA5E]=8'h43; rom['hA5F]=8'hBC;
    rom['hA60]=8'h43; rom['hA61]=8'hC8; rom['hA62]=8'h43; rom['hA63]=8'hC9;
    rom['hA64]=8'h43; rom['hA65]=8'hD5; rom['hA66]=8'h43; rom['hA67]=8'hE9;
    rom['hA68]=8'h43; rom['hA69]=8'hED; rom['hA6A]=8'h43; rom['hA6B]=8'hF9;
    rom['hA6C]=8'h44; rom['hA6D]=8'h05; rom['hA6E]=8'h44; rom['hA6F]=8'h0B;
    rom['hA70]=8'h44; rom['hA71]=8'h0D; rom['hA72]=8'h44; rom['hA73]=8'h0E;
    rom['hA74]=8'h44; rom['hA75]=8'h16; rom['hA76]=8'h44; rom['hA77]=8'h2A;
    rom['hA78]=8'h44; rom['hA79]=8'h2E; rom['hA7A]=8'h44; rom['hA7B]=8'h34;
    rom['hA7C]=8'h44; rom['hA7D]=8'h3A; rom['hA7E]=8'h44; rom['hA7F]=8'h40;
    rom['hA80]=8'h44; rom['hA81]=8'h45; rom['hA82]=8'h44; rom['hA83]=8'h49;
    rom['hA84]=8'h44; rom['hA85]=8'h4F; rom['hA86]=8'h44; rom['hA87]=8'h5F;
    rom['hA88]=8'h44; rom['hA89]=8'h6D; rom['hA8A]=8'h44; rom['hA8B]=8'h71;
    rom['hA8C]=8'h44; rom['hA8D]=8'h77; rom['hA8E]=8'h44; rom['hA8F]=8'h81;
    rom['hA90]=8'h44; rom['hA91]=8'h87; rom['hA92]=8'h44; rom['hA93]=8'h8F;
    rom['hA94]=8'h44; rom['hA95]=8'h95; rom['hA96]=8'h44; rom['hA97]=8'h99;
    rom['hA98]=8'h44; rom['hA99]=8'h9A; rom['hA9A]=8'h44; rom['hA9B]=8'hAA;
    rom['hA9C]=8'h44; rom['hA9D]=8'hC2; rom['hA9E]=8'h44; rom['hA9F]=8'hD9;
    rom['hAA0]=8'h44; rom['hAA1]=8'hDF; rom['hAA2]=8'h44; rom['hAA3]=8'hE3;
    rom['hAA4]=8'h44; rom['hAA5]=8'hE9; rom['hAA6]=8'h44; rom['hAA7]=8'hED;
    rom['hAA8]=8'h44; rom['hAA9]=8'hF1; rom['hAAA]=8'h44; rom['hAAB]=8'hF5;
    rom['hAAC]=8'h44; rom['hAAD]=8'hFB; rom['hAAE]=8'h45; rom['hAAF]=8'h05;
    rom['hAB0]=8'h45; rom['hAB1]=8'h0B; rom['hAB2]=8'h45; rom['hAB3]=8'h0F;
    rom['hAB4]=8'h45; rom['hAB5]=8'h10; rom['hAB6]=8'h45; rom['hAB7]=8'h14;
    rom['hAB8]=8'h45; rom['hAB9]=8'h18; rom['hABA]=8'h45; rom['hABB]=8'h1C;
    rom['hABC]=8'h45; rom['hABD]=8'h1D; rom['hABE]=8'h45; rom['hABF]=8'h2D;
    rom['hAC0]=8'h45; rom['hAC1]=8'h33; rom['hAC2]=8'h45; rom['hAC3]=8'h37;
    rom['hAC4]=8'h45; rom['hAC5]=8'h3D; rom['hAC6]=8'h45; rom['hAC7]=8'h41;
    rom['hAC8]=8'h45; rom['hAC9]=8'h65; rom['hACA]=8'h45; rom['hACB]=8'h69;
    rom['hACC]=8'h45; rom['hACD]=8'h6F; rom['hACE]=8'h45; rom['hACF]=8'h81;
    rom['hAD0]=8'h45; rom['hAD1]=8'h87; rom['hAD2]=8'h45; rom['hAD3]=8'h8B;
    rom['hAD4]=8'h45; rom['hAD5]=8'h8F; rom['hAD6]=8'h45; rom['hAD7]=8'h93;
    rom['hAD8]=8'h45; rom['hAD9]=8'hA1; rom['hADA]=8'h45; rom['hADB]=8'hA5;
    rom['hADC]=8'h45; rom['hADD]=8'hA6; rom['hADE]=8'h45; rom['hADF]=8'hB8;
    rom['hAE0]=8'h45; rom['hAE1]=8'hBE; rom['hAE2]=8'h45; rom['hAE3]=8'hC2;
    rom['hAE4]=8'h45; rom['hAE5]=8'hD0; rom['hAE6]=8'h45; rom['hAE7]=8'hD4;
    rom['hAE8]=8'h45; rom['hAE9]=8'hD5; rom['hAEA]=8'h45; rom['hAEB]=8'hD9;
    rom['hAEC]=8'h45; rom['hAED]=8'hEB; rom['hAEE]=8'h45; rom['hAEF]=8'hFD;
    rom['hAF0]=8'h46; rom['hAF1]=8'h03; rom['hAF2]=8'h46; rom['hAF3]=8'h07;
    rom['hAF4]=8'h46; rom['hAF5]=8'h0D; rom['hAF6]=8'h46; rom['hAF7]=8'h11;
    rom['hAF8]=8'h46; rom['hAF9]=8'h12; rom['hAFA]=8'h46; rom['hAFB]=8'h16;
    rom['hAFC]=8'h46; rom['hAFD]=8'h17; rom['hAFE]=8'h46; rom['hAFF]=8'h27;
    rom['hB00]=8'hA9; rom['hB01]=8'hF8; rom['hB02]=8'hB9; rom['hB03]=8'h12;
    rom['hB04]=8'h08; rom['hB05]=8'hA8; rom['hB06]=8'hF8; rom['hB07]=8'hB8;
    rom['hB08]=8'h29; rom['hB09]=8'hA0; rom['hB0A]=8'hE0; rom['hB0B]=8'hA9;
    rom['hB0C]=8'hF8; rom['hB0D]=8'hB9; rom['hB0E]=8'h29; rom['hB0F]=8'hA1;
    rom['hB10]=8'hE0; rom['hB11]=8'hC0; rom['hB12]=8'hA9; rom['hB13]=8'hF8;
    rom['hB14]=8'hB9; rom['hB15]=8'h12; rom['hB16]=8'h1A; rom['hB17]=8'hA8;
    rom['hB18]=8'hF8; rom['hB19]=8'hB8; rom['hB1A]=8'h29; rom['hB1B]=8'hA2;
    rom['hB1C]=8'hE0; rom['hB1D]=8'hA9; rom['hB1E]=8'hF8; rom['hB1F]=8'hB9;
    rom['hB20]=8'h29; rom['hB21]=8'hA3; rom['hB22]=8'hE0; rom['hB23]=8'hC0;
    rom['hB24]=8'hA9; rom['hB25]=8'hF8; rom['hB26]=8'hB9; rom['hB27]=8'h12;
    rom['hB28]=8'h2C; rom['hB29]=8'hA8; rom['hB2A]=8'hF8; rom['hB2B]=8'hB8;
    rom['hB2C]=8'h29; rom['hB2D]=8'hA4; rom['hB2E]=8'hE0; rom['hB2F]=8'hA9;
    rom['hB30]=8'hF8; rom['hB31]=8'hB9; rom['hB32]=8'h29; rom['hB33]=8'hA5;
    rom['hB34]=8'hE0; rom['hB35]=8'hC0; rom['hB36]=8'h29; rom['hB37]=8'hE9;
    rom['hB38]=8'hB1; rom['hB39]=8'h69; rom['hB3A]=8'h29; rom['hB3B]=8'hE9;
    rom['hB3C]=8'hB0; rom['hB3D]=8'h69; rom['hB3E]=8'hA9; rom['hB3F]=8'h1C;
    rom['hB40]=8'h42; rom['hB41]=8'h68; rom['hB42]=8'hC0; rom['hB43]=8'h29;
    rom['hB44]=8'hE9; rom['hB45]=8'hB3; rom['hB46]=8'h69; rom['hB47]=8'h29;
    rom['hB48]=8'hE9; rom['hB49]=8'hB2; rom['hB4A]=8'h69; rom['hB4B]=8'hA9;
    rom['hB4C]=8'h1C; rom['hB4D]=8'h4F; rom['hB4E]=8'h68; rom['hB4F]=8'hC0;
    rom['hB50]=8'h29; rom['hB51]=8'hE9; rom['hB52]=8'hB5; rom['hB53]=8'h69;
    rom['hB54]=8'h29; rom['hB55]=8'hE9; rom['hB56]=8'hB4; rom['hB57]=8'h69;
    rom['hB58]=8'hA9; rom['hB59]=8'h1C; rom['hB5A]=8'h5C; rom['hB5B]=8'h68;
    rom['hB5C]=8'hC0; rom['hB5D]=8'hA0; rom['hB5E]=8'hBC; rom['hB5F]=8'hA1;
    rom['hB60]=8'hBD; rom['hB61]=8'h2D; rom['hB62]=8'hE9; rom['hB63]=8'h2E;
    rom['hB64]=8'h00; rom['hB65]=8'h2F; rom['hB66]=8'hE1; rom['hB67]=8'h6D;
    rom['hB68]=8'h2D; rom['hB69]=8'hE9; rom['hB6A]=8'h2E; rom['hB6B]=8'h40;
    rom['hB6C]=8'h2F; rom['hB6D]=8'hE1; rom['hB6E]=8'h6D; rom['hB6F]=8'h2D;
    rom['hB70]=8'hE9; rom['hB71]=8'hB1; rom['hB72]=8'h6D; rom['hB73]=8'h2D;
    rom['hB74]=8'hE9; rom['hB75]=8'hB0; rom['hB76]=8'h5F; rom['hB77]=8'hFE;
    rom['hB78]=8'hAC; rom['hB79]=8'hB0; rom['hB7A]=8'hAD; rom['hB7B]=8'hF8;
    rom['hB7C]=8'hF8; rom['hB7D]=8'hF8; rom['hB7E]=8'hB1; rom['hB7F]=8'h48;
    rom['hB80]=8'h5B; rom['hB81]=8'h21; rom['hB82]=8'hE9; rom['hB83]=8'h2E;
    rom['hB84]=8'h00; rom['hB85]=8'h2F; rom['hB86]=8'hE1; rom['hB87]=8'h61;
    rom['hB88]=8'h21; rom['hB89]=8'hE9; rom['hB8A]=8'h2E; rom['hB8B]=8'h40;
    rom['hB8C]=8'h2F; rom['hB8D]=8'hE1; rom['hB8E]=8'h61; rom['hB8F]=8'h21;
    rom['hB90]=8'hE9; rom['hB91]=8'hBD; rom['hB92]=8'h61; rom['hB93]=8'h21;
    rom['hB94]=8'hE9; rom['hB95]=8'hBC; rom['hB96]=8'h2D; rom['hB97]=8'hA3;
    rom['hB98]=8'hE3; rom['hB99]=8'hA2; rom['hB9A]=8'hE3; rom['hB9B]=8'hA1;
    rom['hB9C]=8'hF8; rom['hB9D]=8'hF8; rom['hB9E]=8'hF8; rom['hB9F]=8'hB1;
    rom['hBA0]=8'hC0; rom['hBA1]=8'h21; rom['hBA2]=8'hA3; rom['hBA3]=8'hE3;
    rom['hBA4]=8'hA2; rom['hBA5]=8'hE3; rom['hBA6]=8'hC0; rom['hBA7]=8'h2D;
    rom['hBA8]=8'hAF; rom['hBA9]=8'hE3; rom['hBAA]=8'hAE; rom['hBAB]=8'hE3;
    rom['hBAC]=8'hC0; rom['hBAD]=8'h2C; rom['hBAE]=8'hFE; rom['hBAF]=8'h2E;
    rom['hBB0]=8'h32; rom['hBB1]=8'h5B; rom['hBB2]=8'hA7; rom['hBB3]=8'h6D;
    rom['hBB4]=8'h2E; rom['hBB5]=8'hC0; rom['hBB6]=8'h5B; rom['hBB7]=8'hA7;
    rom['hBB8]=8'hC0; rom['hBB9]=8'h2E; rom['hBBA]=8'h00; rom['hBBB]=8'h2F;
    rom['hBBC]=8'hA3; rom['hBBD]=8'hE1; rom['hBBE]=8'h2E; rom['hBBF]=8'h40;
    rom['hBC0]=8'h2F; rom['hBC1]=8'hA2; rom['hBC2]=8'hE1; rom['hBC3]=8'hC0;
    rom['hBC4]=8'h5B; rom['hBC5]=8'h00; rom['hBC6]=8'h5B; rom['hBC7]=8'h12;
    rom['hBC8]=8'h22; rom['hBC9]=8'h30; rom['hBCA]=8'h57; rom['hBCB]=8'h76;
    rom['hBCC]=8'h5C; rom['hBCD]=8'h37; rom['hBCE]=8'h1C; rom['hBCF]=8'hCC;
    rom['hBD0]=8'h5D; rom['hBD1]=8'h3C; rom['hBD2]=8'h14; rom['hBD3]=8'hDA;
    rom['hBD4]=8'h5C; rom['hBD5]=8'hAC; rom['hBD6]=8'h5C; rom['hBD7]=8'hB0;
    rom['hBD8]=8'h4B; rom['hBD9]=8'hFE; rom['hBDA]=8'h2E; rom['hBDB]=8'h08;
    rom['hBDC]=8'h5D; rom['hBDD]=8'h27; rom['hBDE]=8'h14; rom['hBDF]=8'hE2;
    rom['hBE0]=8'h4B; rom['hBE1]=8'hF6; rom['hBE2]=8'h22; rom['hBE3]=8'h30;
    rom['hBE4]=8'h58; rom['hBE5]=8'h7C; rom['hBE6]=8'h1C; rom['hBE7]=8'hEA;
    rom['hBE8]=8'h4B; rom['hBE9]=8'hCC; rom['hBEA]=8'h58; rom['hBEB]=8'h6B;
    rom['hBEC]=8'h22; rom['hBED]=8'h08; rom['hBEE]=8'h5C; rom['hBEF]=8'h5F;
    rom['hBF0]=8'h5C; rom['hBF1]=8'h98; rom['hBF2]=8'h5C; rom['hBF3]=8'h5F;
    rom['hBF4]=8'h4B; rom['hBF5]=8'hCC; rom['hBF6]=8'h5C; rom['hBF7]=8'h5F;
    rom['hBF8]=8'h5B; rom['hBF9]=8'h81; rom['hBFA]=8'h58; rom['hBFB]=8'h5B;
    rom['hBFC]=8'h4B; rom['hBFD]=8'hCC; rom['hBFE]=8'h22; rom['hBFF]=8'h00;
    rom['hC00]=8'h5B; rom['hC01]=8'h81; rom['hC02]=8'h22; rom['hC03]=8'h30;
    rom['hC04]=8'h57; rom['hC05]=8'h6C; rom['hC06]=8'h5B; rom['hC07]=8'h43;
    rom['hC08]=8'h4B; rom['hC09]=8'h36; rom['hC0A]=8'h5B; rom['hC0B]=8'h12;
    rom['hC0C]=8'h5B; rom['hC0D]=8'h5D; rom['hC0E]=8'h5D; rom['hC0F]=8'h34;
    rom['hC10]=8'h14; rom['hC11]=8'h16; rom['hC12]=8'h5C; rom['hC13]=8'h5F;
    rom['hC14]=8'h4C; rom['hC15]=8'h0C; rom['hC16]=8'h4B; rom['hC17]=8'h43;
    rom['hC18]=8'h5B; rom['hC19]=8'h5D; rom['hC1A]=8'h5C; rom['hC1B]=8'hF0;
    rom['hC1C]=8'h1C; rom['hC1D]=8'h1F; rom['hC1E]=8'hC1; rom['hC1F]=8'h5B;
    rom['hC20]=8'h24; rom['hC21]=8'h5D; rom['hC22]=8'h1B; rom['hC23]=8'hA3;
    rom['hC24]=8'hB4; rom['hC25]=8'h5B; rom['hC26]=8'h5D; rom['hC27]=8'h5C;
    rom['hC28]=8'hF0; rom['hC29]=8'h14; rom['hC2A]=8'h31; rom['hC2B]=8'h5D;
    rom['hC2C]=8'h1B; rom['hC2D]=8'hA4; rom['hC2E]=8'hB2; rom['hC2F]=8'h4B;
    rom['hC30]=8'h50; rom['hC31]=8'hF0; rom['hC32]=8'hB2; rom['hC33]=8'hA4;
    rom['hC34]=8'hB3; rom['hC35]=8'h4B; rom['hC36]=8'h50; rom['hC37]=8'h2C;
    rom['hC38]=8'h0C; rom['hC39]=8'h19; rom['hC3A]=8'h39; rom['hC3B]=8'h2E;
    rom['hC3C]=8'h0C; rom['hC3D]=8'h7F; rom['hC3E]=8'h3D; rom['hC3F]=8'h19;
    rom['hC40]=8'h44; rom['hC41]=8'hF1; rom['hC42]=8'h4C; rom['hC43]=8'h47;
    rom['hC44]=8'hFA; rom['hC45]=8'h00; rom['hC46]=8'h00; rom['hC47]=8'hF6;
    rom['hC48]=8'h00; rom['hC49]=8'h7D; rom['hC4A]=8'h3F; rom['hC4B]=8'hB3;
    rom['hC4C]=8'h2C; rom['hC4D]=8'h0C; rom['hC4E]=8'h19; rom['hC4F]=8'h53;
    rom['hC50]=8'hF1; rom['hC51]=8'h4C; rom['hC52]=8'h56; rom['hC53]=8'hFA;
    rom['hC54]=8'h00; rom['hC55]=8'h00; rom['hC56]=8'hF6; rom['hC57]=8'h00;
    rom['hC58]=8'h7D; rom['hC59]=8'h4E; rom['hC5A]=8'hB2; rom['hC5B]=8'h19;
    rom['hC5C]=8'h5E; rom['hC5D]=8'hC1; rom['hC5E]=8'hC0; rom['hC5F]=8'h2E;
    rom['hC60]=8'hC0; rom['hC61]=8'h2F; rom['hC62]=8'h2C; rom['hC63]=8'h0B;
    rom['hC64]=8'hA3; rom['hC65]=8'hF1; rom['hC66]=8'hF5; rom['hC67]=8'h00;
    rom['hC68]=8'h00; rom['hC69]=8'h00; rom['hC6A]=8'h00; rom['hC6B]=8'h00;
    rom['hC6C]=8'hE1; rom['hC6D]=8'hF6; rom['hC6E]=8'h7D; rom['hC6F]=8'h67;
    rom['hC70]=8'h2C; rom['hC71]=8'h0B; rom['hC72]=8'hA2; rom['hC73]=8'hFA;
    rom['hC74]=8'h00; rom['hC75]=8'h00; rom['hC76]=8'hE1; rom['hC77]=8'h2E;
    rom['hC78]=8'h0E; rom['hC79]=8'h7F; rom['hC7A]=8'h79; rom['hC7B]=8'hF6;
    rom['hC7C]=8'h7D; rom['hC7D]=8'h76; rom['hC7E]=8'hC0; rom['hC7F]=8'h2E;
    rom['hC80]=8'hC0; rom['hC81]=8'h2F; rom['hC82]=8'hD1; rom['hC83]=8'hE1;
    rom['hC84]=8'hC0; rom['hC85]=8'h5B; rom['hC86]=8'h00; rom['hC87]=8'h5B;
    rom['hC88]=8'h12; rom['hC89]=8'hA2; rom['hC8A]=8'hB0; rom['hC8B]=8'hA3;
    rom['hC8C]=8'hB1; rom['hC8D]=8'hA0; rom['hC8E]=8'h5C; rom['hC8F]=8'hB4;
    rom['hC90]=8'hA1; rom['hC91]=8'h5C; rom['hC92]=8'hB4; rom['hC93]=8'h5B;
    rom['hC94]=8'h43; rom['hC95]=8'h5B; rom['hC96]=8'h36; rom['hC97]=8'hC0;
    rom['hC98]=8'h5B; rom['hC99]=8'h12; rom['hC9A]=8'h22; rom['hC9B]=8'h20;
    rom['hC9C]=8'h5C; rom['hC9D]=8'h5F; rom['hC9E]=8'h4B; rom['hC9F]=8'h43;
    rom['hCA0]=8'h5B; rom['hCA1]=8'h12; rom['hCA2]=8'h22; rom['hCA3]=8'h0D;
    rom['hCA4]=8'h5C; rom['hCA5]=8'h5F; rom['hCA6]=8'h22; rom['hCA7]=8'h0A;
    rom['hCA8]=8'h5C; rom['hCA9]=8'h5F; rom['hCAA]=8'h4B; rom['hCAB]=8'h43;
    rom['hCAC]=8'h22; rom['hCAD]=8'h0D; rom['hCAE]=8'h4C; rom['hCAF]=8'h5F;
    rom['hCB0]=8'h22; rom['hCB1]=8'h0A; rom['hCB2]=8'h4C; rom['hCB3]=8'h5F;
    rom['hCB4]=8'h22; rom['hCB5]=8'h30; rom['hCB6]=8'hF1; rom['hCB7]=8'hFB;
    rom['hCB8]=8'h1A; rom['hCB9]=8'hBC; rom['hCBA]=8'h62; rom['hCBB]=8'hF2;
    rom['hCBC]=8'hB3; rom['hCBD]=8'h4C; rom['hCBE]=8'h5F; rom['hCBF]=8'hF0;
    rom['hCC0]=8'h63; rom['hCC1]=8'hA3; rom['hCC2]=8'h1C; rom['hCC3]=8'hC9;
    rom['hCC4]=8'h62; rom['hCC5]=8'hA2; rom['hCC6]=8'h1C; rom['hCC7]=8'hC9;
    rom['hCC8]=8'hFA; rom['hCC9]=8'hC0; rom['hCCA]=8'hA3; rom['hCCB]=8'hF8;
    rom['hCCC]=8'hB3; rom['hCCD]=8'h12; rom['hCCE]=8'hD2; rom['hCCF]=8'hA2;
    rom['hCD0]=8'hF8; rom['hCD1]=8'hB2; rom['hCD2]=8'hC0; rom['hCD3]=8'h2E;
    rom['hCD4]=8'h41; rom['hCD5]=8'h5D; rom['hCD6]=8'h27; rom['hCD7]=8'h12;
    rom['hCD8]=8'hDA; rom['hCD9]=8'hC0; rom['hCDA]=8'h2E; rom['hCDB]=8'h5B;
    rom['hCDC]=8'h5D; rom['hCDD]=8'h27; rom['hCDE]=8'h12; rom['hCDF]=8'hE1;
    rom['hCE0]=8'hC1; rom['hCE1]=8'h2E; rom['hCE2]=8'h61; rom['hCE3]=8'h5D;
    rom['hCE4]=8'h27; rom['hCE5]=8'h12; rom['hCE6]=8'hE8; rom['hCE7]=8'hC0;
    rom['hCE8]=8'h2E; rom['hCE9]=8'h7B; rom['hCEA]=8'h5D; rom['hCEB]=8'h27;
    rom['hCEC]=8'h12; rom['hCED]=8'hEF; rom['hCEE]=8'hC1; rom['hCEF]=8'hC0;
    rom['hCF0]=8'h2E; rom['hCF1]=8'h30; rom['hCF2]=8'h5D; rom['hCF3]=8'h27;
    rom['hCF4]=8'h12; rom['hCF5]=8'hF7; rom['hCF6]=8'hC0; rom['hCF7]=8'h2E;
    rom['hCF8]=8'h3A; rom['hCF9]=8'h5D; rom['hCFA]=8'h27; rom['hCFB]=8'h12;
    rom['hCFC]=8'hFE; rom['hCFD]=8'hC1; rom['hCFE]=8'h2E; rom['hCFF]=8'h41;
    rom['hD00]=8'h5D; rom['hD01]=8'h27; rom['hD02]=8'h12; rom['hD03]=8'h05;
    rom['hD04]=8'hC0; rom['hD05]=8'h2E; rom['hD06]=8'h47; rom['hD07]=8'h5D;
    rom['hD08]=8'h27; rom['hD09]=8'h12; rom['hD0A]=8'h0C; rom['hD0B]=8'hC1;
    rom['hD0C]=8'h2E; rom['hD0D]=8'h61; rom['hD0E]=8'h5D; rom['hD0F]=8'h27;
    rom['hD10]=8'h12; rom['hD11]=8'h13; rom['hD12]=8'hC0; rom['hD13]=8'h2E;
    rom['hD14]=8'h67; rom['hD15]=8'h5D; rom['hD16]=8'h27; rom['hD17]=8'h12;
    rom['hD18]=8'h1A; rom['hD19]=8'hC1; rom['hD1A]=8'hC0; rom['hD1B]=8'hF0;
    rom['hD1C]=8'hD3; rom['hD1D]=8'h92; rom['hD1E]=8'h14; rom['hD1F]=8'h24;
    rom['hD20]=8'hF0; rom['hD21]=8'hD9; rom['hD22]=8'h83; rom['hD23]=8'hB3;
    rom['hD24]=8'hF0; rom['hD25]=8'hB2; rom['hD26]=8'hC0; rom['hD27]=8'hF0;
    rom['hD28]=8'hA2; rom['hD29]=8'h9E; rom['hD2A]=8'h14; rom['hD2B]=8'h2D;
    rom['hD2C]=8'hC1; rom['hD2D]=8'hF0; rom['hD2E]=8'hA3; rom['hD2F]=8'h9F;
    rom['hD30]=8'h14; rom['hD31]=8'h33; rom['hD32]=8'hC1; rom['hD33]=8'hC0;
    rom['hD34]=8'hA3; rom['hD35]=8'h1C; rom['hD36]=8'h3B; rom['hD37]=8'hA2;
    rom['hD38]=8'h1C; rom['hD39]=8'h3B; rom['hD3A]=8'hC0; rom['hD3B]=8'hC1;
    rom['hD3C]=8'hA2; rom['hD3D]=8'h1C; rom['hD3E]=8'h49; rom['hD3F]=8'hF1;
    rom['hD40]=8'hDD; rom['hD41]=8'h93; rom['hD42]=8'h14; rom['hD43]=8'h4A;
    rom['hD44]=8'hF1; rom['hD45]=8'hDA; rom['hD46]=8'h93; rom['hD47]=8'h14;
    rom['hD48]=8'h4A; rom['hD49]=8'hC0; rom['hD4A]=8'hC1; rom['hD4B]=8'h5C;
    rom['hD4C]=8'hD3; rom['hD4D]=8'h14; rom['hD4E]=8'h56; rom['hD4F]=8'hA2;
    rom['hD50]=8'hF6; rom['hD51]=8'hF6; rom['hD52]=8'hF1; rom['hD53]=8'hF5;
    rom['hD54]=8'hF5; rom['hD55]=8'hB2; rom['hD56]=8'hC0; rom['hD57]=8'hA0;
    rom['hD58]=8'h5C; rom['hD59]=8'hB4; rom['hD5A]=8'hA1; rom['hD5B]=8'h5C;
    rom['hD5C]=8'hB4; rom['hD5D]=8'h22; rom['hD5E]=8'h3A; rom['hD5F]=8'h5C;
    rom['hD60]=8'h5F; rom['hD61]=8'hF0; rom['hD62]=8'h21; rom['hD63]=8'hE9;
    rom['hD64]=8'h5C; rom['hD65]=8'hB4; rom['hD66]=8'h71; rom['hD67]=8'h61;
    rom['hD68]=8'h22; rom['hD69]=8'h3A; rom['hD6A]=8'h5C; rom['hD6B]=8'h5F;
    rom['hD6C]=8'h21; rom['hD6D]=8'hEC; rom['hD6E]=8'hB2; rom['hD6F]=8'hED;
    rom['hD70]=8'hB3; rom['hD71]=8'h5C; rom['hD72]=8'h85; rom['hD73]=8'h21;
    rom['hD74]=8'hEE; rom['hD75]=8'hB2; rom['hD76]=8'hEF; rom['hD77]=8'hB3;
    rom['hD78]=8'h5C; rom['hD79]=8'h85; rom['hD7A]=8'h4C; rom['hD7B]=8'hA0;
    rom['hD7C]=8'hFF; rom['hD7D]=8'hFF; rom['hD7E]=8'hFF; rom['hD7F]=8'hFF;
    rom['hD80]=8'hFF; rom['hD81]=8'hFF; rom['hD82]=8'hFF; rom['hD83]=8'hFF;
    rom['hD84]=8'hFF; rom['hD85]=8'hFF; rom['hD86]=8'hFF; rom['hD87]=8'hFF;
    rom['hD88]=8'hFF; rom['hD89]=8'hFF; rom['hD8A]=8'hFF; rom['hD8B]=8'hFF;
    rom['hD8C]=8'hFF; rom['hD8D]=8'hFF; rom['hD8E]=8'hFF; rom['hD8F]=8'hFF;
    rom['hD90]=8'hFF; rom['hD91]=8'hFF; rom['hD92]=8'hFF; rom['hD93]=8'hFF;
    rom['hD94]=8'hFF; rom['hD95]=8'hFF; rom['hD96]=8'hFF; rom['hD97]=8'hFF;
    rom['hD98]=8'hFF; rom['hD99]=8'hFF; rom['hD9A]=8'hFF; rom['hD9B]=8'hFF;
    rom['hD9C]=8'hFF; rom['hD9D]=8'hFF; rom['hD9E]=8'hFF; rom['hD9F]=8'hFF;
    rom['hDA0]=8'hFF; rom['hDA1]=8'hFF; rom['hDA2]=8'hFF; rom['hDA3]=8'hFF;
    rom['hDA4]=8'hFF; rom['hDA5]=8'hFF; rom['hDA6]=8'hFF; rom['hDA7]=8'hFF;
    rom['hDA8]=8'hFF; rom['hDA9]=8'hFF; rom['hDAA]=8'hFF; rom['hDAB]=8'hFF;
    rom['hDAC]=8'hFF; rom['hDAD]=8'hFF; rom['hDAE]=8'hFF; rom['hDAF]=8'hFF;
    rom['hDB0]=8'hFF; rom['hDB1]=8'hFF; rom['hDB2]=8'hFF; rom['hDB3]=8'hFF;
    rom['hDB4]=8'hFF; rom['hDB5]=8'hFF; rom['hDB6]=8'hFF; rom['hDB7]=8'hFF;
    rom['hDB8]=8'hFF; rom['hDB9]=8'hFF; rom['hDBA]=8'hFF; rom['hDBB]=8'hFF;
    rom['hDBC]=8'hFF; rom['hDBD]=8'hFF; rom['hDBE]=8'hFF; rom['hDBF]=8'hFF;
    rom['hDC0]=8'hFF; rom['hDC1]=8'hFF; rom['hDC2]=8'hFF; rom['hDC3]=8'hFF;
    rom['hDC4]=8'hFF; rom['hDC5]=8'hFF; rom['hDC6]=8'hFF; rom['hDC7]=8'hFF;
    rom['hDC8]=8'hFF; rom['hDC9]=8'hFF; rom['hDCA]=8'hFF; rom['hDCB]=8'hFF;
    rom['hDCC]=8'hFF; rom['hDCD]=8'hFF; rom['hDCE]=8'hFF; rom['hDCF]=8'hFF;
    rom['hDD0]=8'hFF; rom['hDD1]=8'hFF; rom['hDD2]=8'hFF; rom['hDD3]=8'hFF;
    rom['hDD4]=8'hFF; rom['hDD5]=8'hFF; rom['hDD6]=8'hFF; rom['hDD7]=8'hFF;
    rom['hDD8]=8'hFF; rom['hDD9]=8'hFF; rom['hDDA]=8'hFF; rom['hDDB]=8'hFF;
    rom['hDDC]=8'hFF; rom['hDDD]=8'hFF; rom['hDDE]=8'hFF; rom['hDDF]=8'hFF;
    rom['hDE0]=8'hFF; rom['hDE1]=8'hFF; rom['hDE2]=8'hFF; rom['hDE3]=8'hFF;
    rom['hDE4]=8'hFF; rom['hDE5]=8'hFF; rom['hDE6]=8'hFF; rom['hDE7]=8'hFF;
    rom['hDE8]=8'hFF; rom['hDE9]=8'hFF; rom['hDEA]=8'hFF; rom['hDEB]=8'hFF;
    rom['hDEC]=8'hFF; rom['hDED]=8'hFF; rom['hDEE]=8'hFF; rom['hDEF]=8'hFF;
    rom['hDF0]=8'hFF; rom['hDF1]=8'hFF; rom['hDF2]=8'hFF; rom['hDF3]=8'hFF;
    rom['hDF4]=8'hFF; rom['hDF5]=8'hFF; rom['hDF6]=8'hFF; rom['hDF7]=8'hFF;
    rom['hDF8]=8'hFF; rom['hDF9]=8'hFF; rom['hDFA]=8'hFF; rom['hDFB]=8'hFF;
    rom['hDFC]=8'hFF; rom['hDFD]=8'hFF; rom['hDFE]=8'hFF; rom['hDFF]=8'hFF;
    rom['hE00]=8'h5B; rom['hE01]=8'h00; rom['hE02]=8'h5B; rom['hE03]=8'h12;
    rom['hE04]=8'h32; rom['hE05]=8'hA2; rom['hE06]=8'h1C; rom['hE07]=8'h0B;
    rom['hE08]=8'hA3; rom['hE09]=8'h14; rom['hE0A]=8'h12; rom['hE0B]=8'h5C;
    rom['hE0C]=8'h5F; rom['hE0D]=8'h71; rom['hE0E]=8'h04; rom['hE0F]=8'h60;
    rom['hE10]=8'h4E; rom['hE11]=8'h04; rom['hE12]=8'h5B; rom['hE13]=8'h43;
    rom['hE14]=8'h4B; rom['hE15]=8'h36; rom['hE16]=8'hA5; rom['hE17]=8'hB4;
    rom['hE18]=8'hA6; rom['hE19]=8'hB5; rom['hE1A]=8'hA7; rom['hE1B]=8'hB6;
    rom['hE1C]=8'hF0; rom['hE1D]=8'hB7; rom['hE1E]=8'hC0; rom['hE1F]=8'h0D;
    rom['hE20]=8'h49; rom['hE21]=8'h6E; rom['hE22]=8'h74; rom['hE23]=8'h65;
    rom['hE24]=8'h6C; rom['hE25]=8'h20; rom['hE26]=8'h4D; rom['hE27]=8'h43;
    rom['hE28]=8'h53; rom['hE29]=8'h2D; rom['hE2A]=8'h34; rom['hE2B]=8'h20;
    rom['hE2C]=8'h28; rom['hE2D]=8'h34; rom['hE2E]=8'h30; rom['hE2F]=8'h30;
    rom['hE30]=8'h34; rom['hE31]=8'h29; rom['hE32]=8'h20; rom['hE33]=8'h54;
    rom['hE34]=8'h69; rom['hE35]=8'h6E; rom['hE36]=8'h79; rom['hE37]=8'h20;
    rom['hE38]=8'h4D; rom['hE39]=8'h6F; rom['hE3A]=8'h6E; rom['hE3B]=8'h69;
    rom['hE3C]=8'h74; rom['hE3D]=8'h6F; rom['hE3E]=8'h72; rom['hE3F]=8'h0D;
    rom['hE40]=8'h0A; rom['hE41]=8'h00; rom['hE42]=8'h1B; rom['hE43]=8'h40;
    rom['hE44]=8'h1F; rom['hE45]=8'h02; rom['hE46]=8'h00; rom['hE47]=8'h3F;
    rom['hE48]=8'h0D; rom['hE49]=8'h0A; rom['hE4A]=8'h00; rom['hE4B]=8'h3F;
    rom['hE4C]=8'h4D; rom['hE4D]=8'h45; rom['hE4E]=8'h4D; rom['hE4F]=8'h53;
    rom['hE50]=8'h50; rom['hE51]=8'h41; rom['hE52]=8'h43; rom['hE53]=8'h45;
    rom['hE54]=8'h0D; rom['hE55]=8'h0A; rom['hE56]=8'h00; rom['hE57]=8'h3F;
    rom['hE58]=8'h4C; rom['hE59]=8'h4F; rom['hE5A]=8'h41; rom['hE5B]=8'h44;
    rom['hE5C]=8'h20; rom['hE5D]=8'h45; rom['hE5E]=8'h52; rom['hE5F]=8'h52;
    rom['hE60]=8'h4F; rom['hE61]=8'h52; rom['hE62]=8'h0D; rom['hE63]=8'h0A;
    rom['hE64]=8'h00; rom['hE65]=8'h0D; rom['hE66]=8'h0A; rom['hE67]=8'h38;
    rom['hE68]=8'h30; rom['hE69]=8'h38; rom['hE6A]=8'h30; rom['hE6B]=8'h20;
    rom['hE6C]=8'h45; rom['hE6D]=8'h6D; rom['hE6E]=8'h75; rom['hE6F]=8'h6C;
    rom['hE70]=8'h61; rom['hE71]=8'h74; rom['hE72]=8'h6F; rom['hE73]=8'h72;
    rom['hE74]=8'h20; rom['hE75]=8'h6F; rom['hE76]=8'h6E; rom['hE77]=8'h20;
    rom['hE78]=8'h34; rom['hE79]=8'h30; rom['hE7A]=8'h30; rom['hE7B]=8'h34;
    rom['hE7C]=8'h20; rom['hE7D]=8'h56; rom['hE7E]=8'h65; rom['hE7F]=8'h72;
    rom['hE80]=8'h20; rom['hE81]=8'h32; rom['hE82]=8'h2E; rom['hE83]=8'h30;
    rom['hE84]=8'h0D; rom['hE85]=8'h0A; rom['hE86]=8'h00; rom['hE87]=8'h41;
    rom['hE88]=8'h20; rom['hE89]=8'h20; rom['hE8A]=8'h53; rom['hE8B]=8'h5A;
    rom['hE8C]=8'h43; rom['hE8D]=8'h20; rom['hE8E]=8'h20; rom['hE8F]=8'h42;
    rom['hE90]=8'h43; rom['hE91]=8'h20; rom['hE92]=8'h20; rom['hE93]=8'h20;
    rom['hE94]=8'h44; rom['hE95]=8'h45; rom['hE96]=8'h20; rom['hE97]=8'h20;
    rom['hE98]=8'h20; rom['hE99]=8'h48; rom['hE9A]=8'h4C; rom['hE9B]=8'h20;
    rom['hE9C]=8'h20; rom['hE9D]=8'h20; rom['hE9E]=8'h53; rom['hE9F]=8'h50;
    rom['hEA0]=8'h20; rom['hEA1]=8'h20; rom['hEA2]=8'h20; rom['hEA3]=8'h50;
    rom['hEA4]=8'h43; rom['hEA5]=8'h20; rom['hEA6]=8'h28; rom['hEA7]=8'h2B;
    rom['hEA8]=8'h30; rom['hEA9]=8'h20; rom['hEAA]=8'h2B; rom['hEAB]=8'h31;
    rom['hEAC]=8'h20; rom['hEAD]=8'h2B; rom['hEAE]=8'h32; rom['hEAF]=8'h29;
    rom['hEB0]=8'h42; rom['hEB1]=8'h43; rom['hEB2]=8'h29; rom['hEB3]=8'h44;
    rom['hEB4]=8'h45; rom['hEB5]=8'h29; rom['hEB6]=8'h48; rom['hEB7]=8'h4C;
    rom['hEB8]=8'h29; rom['hEB9]=8'h53; rom['hEBA]=8'h50; rom['hEBB]=8'h20;
    rom['hEBC]=8'h2B; rom['hEBD]=8'h31; rom['hEBE]=8'h29; rom['hEBF]=8'h0D;
    rom['hEC0]=8'h0A; rom['hEC1]=8'h00; rom['hEC2]=8'h0D; rom['hEC3]=8'h0A;
    rom['hEC4]=8'h53; rom['hEC5]=8'h54; rom['hEC6]=8'h4F; rom['hEC7]=8'h50;
    rom['hEC8]=8'h0D; rom['hEC9]=8'h0A; rom['hECA]=8'h00; rom['hECB]=8'h0D;
    rom['hECC]=8'h0A; rom['hECD]=8'h48; rom['hECE]=8'h4C; rom['hECF]=8'h54;
    rom['hED0]=8'h0D; rom['hED1]=8'h0A; rom['hED2]=8'h00; rom['hED3]=8'h32;
    rom['hED4]=8'hC0; rom['hED5]=8'h00; rom['hED6]=8'h00; rom['hED7]=8'h00;
    rom['hED8]=8'h00; rom['hED9]=8'h00; rom['hEDA]=8'h00; rom['hEDB]=8'h00;
    rom['hEDC]=8'h00; rom['hEDD]=8'h00; rom['hEDE]=8'h00; rom['hEDF]=8'h00;
    rom['hEE0]=8'h00; rom['hEE1]=8'h00; rom['hEE2]=8'h00; rom['hEE3]=8'h00;
    rom['hEE4]=8'h00; rom['hEE5]=8'h00; rom['hEE6]=8'h00; rom['hEE7]=8'h00;
    rom['hEE8]=8'h00; rom['hEE9]=8'h00; rom['hEEA]=8'h00; rom['hEEB]=8'h00;
    rom['hEEC]=8'h00; rom['hEED]=8'h00; rom['hEEE]=8'h00; rom['hEEF]=8'h00;
    rom['hEF0]=8'h00; rom['hEF1]=8'h00; rom['hEF2]=8'h00; rom['hEF3]=8'h00;
    rom['hEF4]=8'h00; rom['hEF5]=8'h00; rom['hEF6]=8'h00; rom['hEF7]=8'h00;
    rom['hEF8]=8'h00; rom['hEF9]=8'h00; rom['hEFA]=8'h00; rom['hEFB]=8'h00;
    rom['hEFC]=8'h00; rom['hEFD]=8'h00; rom['hEFE]=8'h00; rom['hEFF]=8'h00;
    rom['hF00]=8'h00; rom['hF01]=8'h00; rom['hF02]=8'h00; rom['hF03]=8'h00;
    rom['hF04]=8'h00; rom['hF05]=8'h00; rom['hF06]=8'h00; rom['hF07]=8'h00;
    rom['hF08]=8'h00; rom['hF09]=8'h00; rom['hF0A]=8'h00; rom['hF0B]=8'h00;
    rom['hF0C]=8'h00; rom['hF0D]=8'h00; rom['hF0E]=8'h00; rom['hF0F]=8'h00;
    rom['hF10]=8'h00; rom['hF11]=8'h00; rom['hF12]=8'h00; rom['hF13]=8'h00;
    rom['hF14]=8'h00; rom['hF15]=8'h00; rom['hF16]=8'h00; rom['hF17]=8'h00;
    rom['hF18]=8'h00; rom['hF19]=8'h00; rom['hF1A]=8'h00; rom['hF1B]=8'h00;
    rom['hF1C]=8'h00; rom['hF1D]=8'h00; rom['hF1E]=8'h00; rom['hF1F]=8'h00;
    rom['hF20]=8'h00; rom['hF21]=8'h00; rom['hF22]=8'h00; rom['hF23]=8'h00;
    rom['hF24]=8'h00; rom['hF25]=8'h00; rom['hF26]=8'h00; rom['hF27]=8'h00;
    rom['hF28]=8'h00; rom['hF29]=8'h00; rom['hF2A]=8'h00; rom['hF2B]=8'h00;
    rom['hF2C]=8'h00; rom['hF2D]=8'h00; rom['hF2E]=8'h00; rom['hF2F]=8'h00;
    rom['hF30]=8'h00; rom['hF31]=8'h00; rom['hF32]=8'h00; rom['hF33]=8'h00;
    rom['hF34]=8'h00; rom['hF35]=8'h00; rom['hF36]=8'h00; rom['hF37]=8'h00;
    rom['hF38]=8'h00; rom['hF39]=8'h00; rom['hF3A]=8'h00; rom['hF3B]=8'h00;
    rom['hF3C]=8'h00; rom['hF3D]=8'h00; rom['hF3E]=8'h00; rom['hF3F]=8'h00;
    rom['hF40]=8'h00; rom['hF41]=8'h00; rom['hF42]=8'h00; rom['hF43]=8'h00;
    rom['hF44]=8'h00; rom['hF45]=8'h00; rom['hF46]=8'h00; rom['hF47]=8'h00;
    rom['hF48]=8'h00; rom['hF49]=8'h00; rom['hF4A]=8'h00; rom['hF4B]=8'h00;
    rom['hF4C]=8'h00; rom['hF4D]=8'h00; rom['hF4E]=8'h00; rom['hF4F]=8'h00;
    rom['hF50]=8'h00; rom['hF51]=8'h00; rom['hF52]=8'h00; rom['hF53]=8'h00;
    rom['hF54]=8'h00; rom['hF55]=8'h00; rom['hF56]=8'h00; rom['hF57]=8'h00;
    rom['hF58]=8'h00; rom['hF59]=8'h00; rom['hF5A]=8'h00; rom['hF5B]=8'h00;
    rom['hF5C]=8'h00; rom['hF5D]=8'h00; rom['hF5E]=8'h00; rom['hF5F]=8'h00;
    rom['hF60]=8'h00; rom['hF61]=8'h00; rom['hF62]=8'h00; rom['hF63]=8'h00;
    rom['hF64]=8'h00; rom['hF65]=8'h00; rom['hF66]=8'h00; rom['hF67]=8'h00;
    rom['hF68]=8'h00; rom['hF69]=8'h00; rom['hF6A]=8'h00; rom['hF6B]=8'h00;
    rom['hF6C]=8'h00; rom['hF6D]=8'h00; rom['hF6E]=8'h00; rom['hF6F]=8'h00;
    rom['hF70]=8'h00; rom['hF71]=8'h00; rom['hF72]=8'h00; rom['hF73]=8'h00;
    rom['hF74]=8'h00; rom['hF75]=8'h00; rom['hF76]=8'h00; rom['hF77]=8'h00;
    rom['hF78]=8'h00; rom['hF79]=8'h00; rom['hF7A]=8'h00; rom['hF7B]=8'h00;
    rom['hF7C]=8'h00; rom['hF7D]=8'h00; rom['hF7E]=8'h00; rom['hF7F]=8'h00;
    rom['hF80]=8'h00; rom['hF81]=8'h00; rom['hF82]=8'h00; rom['hF83]=8'h00;
    rom['hF84]=8'h00; rom['hF85]=8'h00; rom['hF86]=8'h00; rom['hF87]=8'h00;
    rom['hF88]=8'h00; rom['hF89]=8'h00; rom['hF8A]=8'h00; rom['hF8B]=8'h00;
    rom['hF8C]=8'h00; rom['hF8D]=8'h00; rom['hF8E]=8'h00; rom['hF8F]=8'h00;
    rom['hF90]=8'h00; rom['hF91]=8'h00; rom['hF92]=8'h00; rom['hF93]=8'h00;
    rom['hF94]=8'h00; rom['hF95]=8'h00; rom['hF96]=8'h00; rom['hF97]=8'h00;
    rom['hF98]=8'h00; rom['hF99]=8'h00; rom['hF9A]=8'h00; rom['hF9B]=8'h00;
    rom['hF9C]=8'h00; rom['hF9D]=8'h00; rom['hF9E]=8'h00; rom['hF9F]=8'h00;
    rom['hFA0]=8'h00; rom['hFA1]=8'h00; rom['hFA2]=8'h00; rom['hFA3]=8'h00;
    rom['hFA4]=8'h00; rom['hFA5]=8'h00; rom['hFA6]=8'h00; rom['hFA7]=8'h00;
    rom['hFA8]=8'h00; rom['hFA9]=8'h00; rom['hFAA]=8'h00; rom['hFAB]=8'h00;
    rom['hFAC]=8'h00; rom['hFAD]=8'h00; rom['hFAE]=8'h00; rom['hFAF]=8'h00;
    rom['hFB0]=8'h00; rom['hFB1]=8'h00; rom['hFB2]=8'h00; rom['hFB3]=8'h00;
    rom['hFB4]=8'h00; rom['hFB5]=8'h00; rom['hFB6]=8'h00; rom['hFB7]=8'h00;
    rom['hFB8]=8'h00; rom['hFB9]=8'h00; rom['hFBA]=8'h00; rom['hFBB]=8'h00;
    rom['hFBC]=8'h00; rom['hFBD]=8'h00; rom['hFBE]=8'h00; rom['hFBF]=8'h00;
    rom['hFC0]=8'h00; rom['hFC1]=8'h00; rom['hFC2]=8'h00; rom['hFC3]=8'h00;
    rom['hFC4]=8'h00; rom['hFC5]=8'h00; rom['hFC6]=8'h00; rom['hFC7]=8'h00;
    rom['hFC8]=8'h00; rom['hFC9]=8'h00; rom['hFCA]=8'h00; rom['hFCB]=8'h00;
    rom['hFCC]=8'h00; rom['hFCD]=8'h00; rom['hFCE]=8'h00; rom['hFCF]=8'h00;
    rom['hFD0]=8'h00; rom['hFD1]=8'h00; rom['hFD2]=8'h00; rom['hFD3]=8'h00;
    rom['hFD4]=8'h00; rom['hFD5]=8'h00; rom['hFD6]=8'h00; rom['hFD7]=8'h00;
    rom['hFD8]=8'h00; rom['hFD9]=8'h00; rom['hFDA]=8'h00; rom['hFDB]=8'h00;
    rom['hFDC]=8'h00; rom['hFDD]=8'h00; rom['hFDE]=8'h00; rom['hFDF]=8'h00;
    rom['hFE0]=8'h00; rom['hFE1]=8'h00; rom['hFE2]=8'h00; rom['hFE3]=8'h00;
    rom['hFE4]=8'h00; rom['hFE5]=8'h00; rom['hFE6]=8'h00; rom['hFE7]=8'h00;
    rom['hFE8]=8'h00; rom['hFE9]=8'h00; rom['hFEA]=8'h00; rom['hFEB]=8'h00;
    rom['hFEC]=8'h00; rom['hFED]=8'h00; rom['hFEE]=8'h00; rom['hFEF]=8'h00;
    rom['hFF0]=8'h00; rom['hFF1]=8'h00; rom['hFF2]=8'h00; rom['hFF3]=8'h00;
    rom['hFF4]=8'h00; rom['hFF5]=8'h00; rom['hFF6]=8'h00; rom['hFF7]=8'h00;
    rom['hFF8]=8'h00; rom['hFF9]=8'h00; rom['hFFA]=8'h00; rom['hFFB]=8'h00;
    rom['hFFC]=8'h00; rom['hFFD]=8'h00; rom['hFFE]=8'h00; rom['hFFF]=8'h00;
    end
endmodule
